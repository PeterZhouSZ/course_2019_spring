module our(clk,reset,read_base,write_base,num_read,read_size_input,read_ready,write_ready,read_data,
			read_enable,write_enable,finish_read,finish_write,read_addr,write_addr,write_size,read_size_output,write_data,done);
    input wire clk;
    input wire reset;
    input wire[63:0] read_base;
	input wire[63:0] write_base;
	input wire[63:0] num_read;
	input wire[63:0] read_size_input;
	input wire[63:0] read_ready;
	input wire[63:0] write_ready;
	input wire[63:0] read_data;
    output wire read_enable;
	output wire write_enable;
	output wire finish_read;
	output wire finish_write;
    output wire done;
	output wire[63:0] read_addr;
	output wire[63:0] write_addr;
	output wire[63:0] write_size;
	output wire[63:0] read_size_output;
    output wire[63:0] write_data;

	reg[63:0] read_cnt;
	reg[63:0] write_cnt;
	reg[63:0] state;
    reg r_read_enable;
	reg r_write_enable;
	reg r_finish_read;
	reg r_finish_write;
    reg r_done;
	reg[63:0] r_read_addr;
	reg[63:0] r_write_addr;
	reg[63:0] r_write_size;
	reg[63:0] r_read_size_output;
    //reg[63:0] r_read_data;
    reg[63:0] r_write_data;
	reg[63:0] tmp[0:10001];
	reg[63:0] ans[0:10001];
	reg[63:0] kernel[0:8];
    assign read_enable=r_read_enable;
	assign write_enable=r_write_enable;
	assign finish_read=r_finish_read;
	assign finish_write=r_finish_write;
	assign read_addr=r_read_addr;
	assign write_addr=r_write_addr;
	assign write_size=r_write_size;
	assign read_size_output=r_read_size_output;
    assign write_data=r_write_data;
    assign done=r_done;




	parameter IDLE = 64'd0;
	parameter READY_READ = 64'd1;
	parameter WAIT_READ = 64'd2;
	parameter DEAL_READ = 64'd3;
	parameter FINISH = 64'd4;
	parameter READY_WRITE = 64'd5;
	parameter WAIT_WRITE = 64'd6;
    parameter DEAL_WRITE = 64'd7;
	parameter SUSPEND = 64'd8;
    parameter LOOP = 64'd9;
    parameter HANDLING = 64'd10;

    always @(posedge reset or posedge clk)
    begin
        if (reset)
        begin
            state<=IDLE;
            read_cnt<=0;
            write_cnt<=0;
            r_read_enable<=0;
            r_write_enable<=0;
            r_finish_read<=0;
            r_finish_write<=0;
            r_read_addr<=0;
            r_write_addr<=0;
            r_write_size<=0;
            r_read_size_output<=0;
            r_done<=0;
			// kernel<={1,2,1,0,0,0,1,2,1};
        end
        else
        begin
            if (state == IDLE)
            begin
                state<=WAIT_READ;
                r_read_addr<=read_base;
                r_read_size_output<=read_size_input;
                r_read_enable<=1;
            end
            else if (state == WAIT_READ)
            begin
                r_finish_read<=0;
                if (read_ready == 1)
                begin
                    tmp[read_cnt[15:0]]<=read_data;
                    state<= DEAL_READ;
                end
            end
            else if (state == DEAL_READ)
            begin
                if (read_cnt + 1 < num_read)
                begin
                    read_cnt<=read_cnt+1;
                    r_read_addr<=r_read_addr+read_size_input;
                    state<=WAIT_READ;
                    r_finish_read<=1;
                end
                else
                begin
                    state<=HANDLING;
                    r_read_enable<=0;
                    r_finish_read<=0;
                end
            end
            else if (state == HANDLING)
            begin
				ans[0]<=tmp[0]*kernel[4]+tmp[1]*kernel[5]+tmp[100]*kernel[7]+tmp[101]*kernel[8];
				ans[1]<=tmp[0]*kernel[3]+tmp[1]*kernel[4]+tmp[2]*kernel[5]+tmp[100]*kernel[6]+tmp[101]*kernel[7]+tmp[102]*kernel[8];
				ans[2]<=tmp[1]*kernel[3]+tmp[2]*kernel[4]+tmp[3]*kernel[5]+tmp[101]*kernel[6]+tmp[102]*kernel[7]+tmp[103]*kernel[8];
				ans[3]<=tmp[2]*kernel[3]+tmp[3]*kernel[4]+tmp[4]*kernel[5]+tmp[102]*kernel[6]+tmp[103]*kernel[7]+tmp[104]*kernel[8];
				ans[4]<=tmp[3]*kernel[3]+tmp[4]*kernel[4]+tmp[5]*kernel[5]+tmp[103]*kernel[6]+tmp[104]*kernel[7]+tmp[105]*kernel[8];
				ans[5]<=tmp[4]*kernel[3]+tmp[5]*kernel[4]+tmp[6]*kernel[5]+tmp[104]*kernel[6]+tmp[105]*kernel[7]+tmp[106]*kernel[8];
				ans[6]<=tmp[5]*kernel[3]+tmp[6]*kernel[4]+tmp[7]*kernel[5]+tmp[105]*kernel[6]+tmp[106]*kernel[7]+tmp[107]*kernel[8];
				ans[7]<=tmp[6]*kernel[3]+tmp[7]*kernel[4]+tmp[8]*kernel[5]+tmp[106]*kernel[6]+tmp[107]*kernel[7]+tmp[108]*kernel[8];
				ans[8]<=tmp[7]*kernel[3]+tmp[8]*kernel[4]+tmp[9]*kernel[5]+tmp[107]*kernel[6]+tmp[108]*kernel[7]+tmp[109]*kernel[8];
				ans[9]<=tmp[8]*kernel[3]+tmp[9]*kernel[4]+tmp[10]*kernel[5]+tmp[108]*kernel[6]+tmp[109]*kernel[7]+tmp[110]*kernel[8];
				ans[10]<=tmp[9]*kernel[3]+tmp[10]*kernel[4]+tmp[11]*kernel[5]+tmp[109]*kernel[6]+tmp[110]*kernel[7]+tmp[111]*kernel[8];
				ans[11]<=tmp[10]*kernel[3]+tmp[11]*kernel[4]+tmp[12]*kernel[5]+tmp[110]*kernel[6]+tmp[111]*kernel[7]+tmp[112]*kernel[8];
				ans[12]<=tmp[11]*kernel[3]+tmp[12]*kernel[4]+tmp[13]*kernel[5]+tmp[111]*kernel[6]+tmp[112]*kernel[7]+tmp[113]*kernel[8];
				ans[13]<=tmp[12]*kernel[3]+tmp[13]*kernel[4]+tmp[14]*kernel[5]+tmp[112]*kernel[6]+tmp[113]*kernel[7]+tmp[114]*kernel[8];
				ans[14]<=tmp[13]*kernel[3]+tmp[14]*kernel[4]+tmp[15]*kernel[5]+tmp[113]*kernel[6]+tmp[114]*kernel[7]+tmp[115]*kernel[8];
				ans[15]<=tmp[14]*kernel[3]+tmp[15]*kernel[4]+tmp[16]*kernel[5]+tmp[114]*kernel[6]+tmp[115]*kernel[7]+tmp[116]*kernel[8];
				ans[16]<=tmp[15]*kernel[3]+tmp[16]*kernel[4]+tmp[17]*kernel[5]+tmp[115]*kernel[6]+tmp[116]*kernel[7]+tmp[117]*kernel[8];
				ans[17]<=tmp[16]*kernel[3]+tmp[17]*kernel[4]+tmp[18]*kernel[5]+tmp[116]*kernel[6]+tmp[117]*kernel[7]+tmp[118]*kernel[8];
				ans[18]<=tmp[17]*kernel[3]+tmp[18]*kernel[4]+tmp[19]*kernel[5]+tmp[117]*kernel[6]+tmp[118]*kernel[7]+tmp[119]*kernel[8];
				ans[19]<=tmp[18]*kernel[3]+tmp[19]*kernel[4]+tmp[20]*kernel[5]+tmp[118]*kernel[6]+tmp[119]*kernel[7]+tmp[120]*kernel[8];
				ans[20]<=tmp[19]*kernel[3]+tmp[20]*kernel[4]+tmp[21]*kernel[5]+tmp[119]*kernel[6]+tmp[120]*kernel[7]+tmp[121]*kernel[8];
				ans[21]<=tmp[20]*kernel[3]+tmp[21]*kernel[4]+tmp[22]*kernel[5]+tmp[120]*kernel[6]+tmp[121]*kernel[7]+tmp[122]*kernel[8];
				ans[22]<=tmp[21]*kernel[3]+tmp[22]*kernel[4]+tmp[23]*kernel[5]+tmp[121]*kernel[6]+tmp[122]*kernel[7]+tmp[123]*kernel[8];
				ans[23]<=tmp[22]*kernel[3]+tmp[23]*kernel[4]+tmp[24]*kernel[5]+tmp[122]*kernel[6]+tmp[123]*kernel[7]+tmp[124]*kernel[8];
				ans[24]<=tmp[23]*kernel[3]+tmp[24]*kernel[4]+tmp[25]*kernel[5]+tmp[123]*kernel[6]+tmp[124]*kernel[7]+tmp[125]*kernel[8];
				ans[25]<=tmp[24]*kernel[3]+tmp[25]*kernel[4]+tmp[26]*kernel[5]+tmp[124]*kernel[6]+tmp[125]*kernel[7]+tmp[126]*kernel[8];
				ans[26]<=tmp[25]*kernel[3]+tmp[26]*kernel[4]+tmp[27]*kernel[5]+tmp[125]*kernel[6]+tmp[126]*kernel[7]+tmp[127]*kernel[8];
				ans[27]<=tmp[26]*kernel[3]+tmp[27]*kernel[4]+tmp[28]*kernel[5]+tmp[126]*kernel[6]+tmp[127]*kernel[7]+tmp[128]*kernel[8];
				ans[28]<=tmp[27]*kernel[3]+tmp[28]*kernel[4]+tmp[29]*kernel[5]+tmp[127]*kernel[6]+tmp[128]*kernel[7]+tmp[129]*kernel[8];
				ans[29]<=tmp[28]*kernel[3]+tmp[29]*kernel[4]+tmp[30]*kernel[5]+tmp[128]*kernel[6]+tmp[129]*kernel[7]+tmp[130]*kernel[8];
				ans[30]<=tmp[29]*kernel[3]+tmp[30]*kernel[4]+tmp[31]*kernel[5]+tmp[129]*kernel[6]+tmp[130]*kernel[7]+tmp[131]*kernel[8];
				ans[31]<=tmp[30]*kernel[3]+tmp[31]*kernel[4]+tmp[32]*kernel[5]+tmp[130]*kernel[6]+tmp[131]*kernel[7]+tmp[132]*kernel[8];
				ans[32]<=tmp[31]*kernel[3]+tmp[32]*kernel[4]+tmp[33]*kernel[5]+tmp[131]*kernel[6]+tmp[132]*kernel[7]+tmp[133]*kernel[8];
				ans[33]<=tmp[32]*kernel[3]+tmp[33]*kernel[4]+tmp[34]*kernel[5]+tmp[132]*kernel[6]+tmp[133]*kernel[7]+tmp[134]*kernel[8];
				ans[34]<=tmp[33]*kernel[3]+tmp[34]*kernel[4]+tmp[35]*kernel[5]+tmp[133]*kernel[6]+tmp[134]*kernel[7]+tmp[135]*kernel[8];
				ans[35]<=tmp[34]*kernel[3]+tmp[35]*kernel[4]+tmp[36]*kernel[5]+tmp[134]*kernel[6]+tmp[135]*kernel[7]+tmp[136]*kernel[8];
				ans[36]<=tmp[35]*kernel[3]+tmp[36]*kernel[4]+tmp[37]*kernel[5]+tmp[135]*kernel[6]+tmp[136]*kernel[7]+tmp[137]*kernel[8];
				ans[37]<=tmp[36]*kernel[3]+tmp[37]*kernel[4]+tmp[38]*kernel[5]+tmp[136]*kernel[6]+tmp[137]*kernel[7]+tmp[138]*kernel[8];
				ans[38]<=tmp[37]*kernel[3]+tmp[38]*kernel[4]+tmp[39]*kernel[5]+tmp[137]*kernel[6]+tmp[138]*kernel[7]+tmp[139]*kernel[8];
				ans[39]<=tmp[38]*kernel[3]+tmp[39]*kernel[4]+tmp[40]*kernel[5]+tmp[138]*kernel[6]+tmp[139]*kernel[7]+tmp[140]*kernel[8];
				ans[40]<=tmp[39]*kernel[3]+tmp[40]*kernel[4]+tmp[41]*kernel[5]+tmp[139]*kernel[6]+tmp[140]*kernel[7]+tmp[141]*kernel[8];
				ans[41]<=tmp[40]*kernel[3]+tmp[41]*kernel[4]+tmp[42]*kernel[5]+tmp[140]*kernel[6]+tmp[141]*kernel[7]+tmp[142]*kernel[8];
				ans[42]<=tmp[41]*kernel[3]+tmp[42]*kernel[4]+tmp[43]*kernel[5]+tmp[141]*kernel[6]+tmp[142]*kernel[7]+tmp[143]*kernel[8];
				ans[43]<=tmp[42]*kernel[3]+tmp[43]*kernel[4]+tmp[44]*kernel[5]+tmp[142]*kernel[6]+tmp[143]*kernel[7]+tmp[144]*kernel[8];
				ans[44]<=tmp[43]*kernel[3]+tmp[44]*kernel[4]+tmp[45]*kernel[5]+tmp[143]*kernel[6]+tmp[144]*kernel[7]+tmp[145]*kernel[8];
				ans[45]<=tmp[44]*kernel[3]+tmp[45]*kernel[4]+tmp[46]*kernel[5]+tmp[144]*kernel[6]+tmp[145]*kernel[7]+tmp[146]*kernel[8];
				ans[46]<=tmp[45]*kernel[3]+tmp[46]*kernel[4]+tmp[47]*kernel[5]+tmp[145]*kernel[6]+tmp[146]*kernel[7]+tmp[147]*kernel[8];
				ans[47]<=tmp[46]*kernel[3]+tmp[47]*kernel[4]+tmp[48]*kernel[5]+tmp[146]*kernel[6]+tmp[147]*kernel[7]+tmp[148]*kernel[8];
				ans[48]<=tmp[47]*kernel[3]+tmp[48]*kernel[4]+tmp[49]*kernel[5]+tmp[147]*kernel[6]+tmp[148]*kernel[7]+tmp[149]*kernel[8];
				ans[49]<=tmp[48]*kernel[3]+tmp[49]*kernel[4]+tmp[50]*kernel[5]+tmp[148]*kernel[6]+tmp[149]*kernel[7]+tmp[150]*kernel[8];
				ans[50]<=tmp[49]*kernel[3]+tmp[50]*kernel[4]+tmp[51]*kernel[5]+tmp[149]*kernel[6]+tmp[150]*kernel[7]+tmp[151]*kernel[8];
				ans[51]<=tmp[50]*kernel[3]+tmp[51]*kernel[4]+tmp[52]*kernel[5]+tmp[150]*kernel[6]+tmp[151]*kernel[7]+tmp[152]*kernel[8];
				ans[52]<=tmp[51]*kernel[3]+tmp[52]*kernel[4]+tmp[53]*kernel[5]+tmp[151]*kernel[6]+tmp[152]*kernel[7]+tmp[153]*kernel[8];
				ans[53]<=tmp[52]*kernel[3]+tmp[53]*kernel[4]+tmp[54]*kernel[5]+tmp[152]*kernel[6]+tmp[153]*kernel[7]+tmp[154]*kernel[8];
				ans[54]<=tmp[53]*kernel[3]+tmp[54]*kernel[4]+tmp[55]*kernel[5]+tmp[153]*kernel[6]+tmp[154]*kernel[7]+tmp[155]*kernel[8];
				ans[55]<=tmp[54]*kernel[3]+tmp[55]*kernel[4]+tmp[56]*kernel[5]+tmp[154]*kernel[6]+tmp[155]*kernel[7]+tmp[156]*kernel[8];
				ans[56]<=tmp[55]*kernel[3]+tmp[56]*kernel[4]+tmp[57]*kernel[5]+tmp[155]*kernel[6]+tmp[156]*kernel[7]+tmp[157]*kernel[8];
				ans[57]<=tmp[56]*kernel[3]+tmp[57]*kernel[4]+tmp[58]*kernel[5]+tmp[156]*kernel[6]+tmp[157]*kernel[7]+tmp[158]*kernel[8];
				ans[58]<=tmp[57]*kernel[3]+tmp[58]*kernel[4]+tmp[59]*kernel[5]+tmp[157]*kernel[6]+tmp[158]*kernel[7]+tmp[159]*kernel[8];
				ans[59]<=tmp[58]*kernel[3]+tmp[59]*kernel[4]+tmp[60]*kernel[5]+tmp[158]*kernel[6]+tmp[159]*kernel[7]+tmp[160]*kernel[8];
				ans[60]<=tmp[59]*kernel[3]+tmp[60]*kernel[4]+tmp[61]*kernel[5]+tmp[159]*kernel[6]+tmp[160]*kernel[7]+tmp[161]*kernel[8];
				ans[61]<=tmp[60]*kernel[3]+tmp[61]*kernel[4]+tmp[62]*kernel[5]+tmp[160]*kernel[6]+tmp[161]*kernel[7]+tmp[162]*kernel[8];
				ans[62]<=tmp[61]*kernel[3]+tmp[62]*kernel[4]+tmp[63]*kernel[5]+tmp[161]*kernel[6]+tmp[162]*kernel[7]+tmp[163]*kernel[8];
				ans[63]<=tmp[62]*kernel[3]+tmp[63]*kernel[4]+tmp[64]*kernel[5]+tmp[162]*kernel[6]+tmp[163]*kernel[7]+tmp[164]*kernel[8];
				ans[64]<=tmp[63]*kernel[3]+tmp[64]*kernel[4]+tmp[65]*kernel[5]+tmp[163]*kernel[6]+tmp[164]*kernel[7]+tmp[165]*kernel[8];
				ans[65]<=tmp[64]*kernel[3]+tmp[65]*kernel[4]+tmp[66]*kernel[5]+tmp[164]*kernel[6]+tmp[165]*kernel[7]+tmp[166]*kernel[8];
				ans[66]<=tmp[65]*kernel[3]+tmp[66]*kernel[4]+tmp[67]*kernel[5]+tmp[165]*kernel[6]+tmp[166]*kernel[7]+tmp[167]*kernel[8];
				ans[67]<=tmp[66]*kernel[3]+tmp[67]*kernel[4]+tmp[68]*kernel[5]+tmp[166]*kernel[6]+tmp[167]*kernel[7]+tmp[168]*kernel[8];
				ans[68]<=tmp[67]*kernel[3]+tmp[68]*kernel[4]+tmp[69]*kernel[5]+tmp[167]*kernel[6]+tmp[168]*kernel[7]+tmp[169]*kernel[8];
				ans[69]<=tmp[68]*kernel[3]+tmp[69]*kernel[4]+tmp[70]*kernel[5]+tmp[168]*kernel[6]+tmp[169]*kernel[7]+tmp[170]*kernel[8];
				ans[70]<=tmp[69]*kernel[3]+tmp[70]*kernel[4]+tmp[71]*kernel[5]+tmp[169]*kernel[6]+tmp[170]*kernel[7]+tmp[171]*kernel[8];
				ans[71]<=tmp[70]*kernel[3]+tmp[71]*kernel[4]+tmp[72]*kernel[5]+tmp[170]*kernel[6]+tmp[171]*kernel[7]+tmp[172]*kernel[8];
				ans[72]<=tmp[71]*kernel[3]+tmp[72]*kernel[4]+tmp[73]*kernel[5]+tmp[171]*kernel[6]+tmp[172]*kernel[7]+tmp[173]*kernel[8];
				ans[73]<=tmp[72]*kernel[3]+tmp[73]*kernel[4]+tmp[74]*kernel[5]+tmp[172]*kernel[6]+tmp[173]*kernel[7]+tmp[174]*kernel[8];
				ans[74]<=tmp[73]*kernel[3]+tmp[74]*kernel[4]+tmp[75]*kernel[5]+tmp[173]*kernel[6]+tmp[174]*kernel[7]+tmp[175]*kernel[8];
				ans[75]<=tmp[74]*kernel[3]+tmp[75]*kernel[4]+tmp[76]*kernel[5]+tmp[174]*kernel[6]+tmp[175]*kernel[7]+tmp[176]*kernel[8];
				ans[76]<=tmp[75]*kernel[3]+tmp[76]*kernel[4]+tmp[77]*kernel[5]+tmp[175]*kernel[6]+tmp[176]*kernel[7]+tmp[177]*kernel[8];
				ans[77]<=tmp[76]*kernel[3]+tmp[77]*kernel[4]+tmp[78]*kernel[5]+tmp[176]*kernel[6]+tmp[177]*kernel[7]+tmp[178]*kernel[8];
				ans[78]<=tmp[77]*kernel[3]+tmp[78]*kernel[4]+tmp[79]*kernel[5]+tmp[177]*kernel[6]+tmp[178]*kernel[7]+tmp[179]*kernel[8];
				ans[79]<=tmp[78]*kernel[3]+tmp[79]*kernel[4]+tmp[80]*kernel[5]+tmp[178]*kernel[6]+tmp[179]*kernel[7]+tmp[180]*kernel[8];
				ans[80]<=tmp[79]*kernel[3]+tmp[80]*kernel[4]+tmp[81]*kernel[5]+tmp[179]*kernel[6]+tmp[180]*kernel[7]+tmp[181]*kernel[8];
				ans[81]<=tmp[80]*kernel[3]+tmp[81]*kernel[4]+tmp[82]*kernel[5]+tmp[180]*kernel[6]+tmp[181]*kernel[7]+tmp[182]*kernel[8];
				ans[82]<=tmp[81]*kernel[3]+tmp[82]*kernel[4]+tmp[83]*kernel[5]+tmp[181]*kernel[6]+tmp[182]*kernel[7]+tmp[183]*kernel[8];
				ans[83]<=tmp[82]*kernel[3]+tmp[83]*kernel[4]+tmp[84]*kernel[5]+tmp[182]*kernel[6]+tmp[183]*kernel[7]+tmp[184]*kernel[8];
				ans[84]<=tmp[83]*kernel[3]+tmp[84]*kernel[4]+tmp[85]*kernel[5]+tmp[183]*kernel[6]+tmp[184]*kernel[7]+tmp[185]*kernel[8];
				ans[85]<=tmp[84]*kernel[3]+tmp[85]*kernel[4]+tmp[86]*kernel[5]+tmp[184]*kernel[6]+tmp[185]*kernel[7]+tmp[186]*kernel[8];
				ans[86]<=tmp[85]*kernel[3]+tmp[86]*kernel[4]+tmp[87]*kernel[5]+tmp[185]*kernel[6]+tmp[186]*kernel[7]+tmp[187]*kernel[8];
				ans[87]<=tmp[86]*kernel[3]+tmp[87]*kernel[4]+tmp[88]*kernel[5]+tmp[186]*kernel[6]+tmp[187]*kernel[7]+tmp[188]*kernel[8];
				ans[88]<=tmp[87]*kernel[3]+tmp[88]*kernel[4]+tmp[89]*kernel[5]+tmp[187]*kernel[6]+tmp[188]*kernel[7]+tmp[189]*kernel[8];
				ans[89]<=tmp[88]*kernel[3]+tmp[89]*kernel[4]+tmp[90]*kernel[5]+tmp[188]*kernel[6]+tmp[189]*kernel[7]+tmp[190]*kernel[8];
				ans[90]<=tmp[89]*kernel[3]+tmp[90]*kernel[4]+tmp[91]*kernel[5]+tmp[189]*kernel[6]+tmp[190]*kernel[7]+tmp[191]*kernel[8];
				ans[91]<=tmp[90]*kernel[3]+tmp[91]*kernel[4]+tmp[92]*kernel[5]+tmp[190]*kernel[6]+tmp[191]*kernel[7]+tmp[192]*kernel[8];
				ans[92]<=tmp[91]*kernel[3]+tmp[92]*kernel[4]+tmp[93]*kernel[5]+tmp[191]*kernel[6]+tmp[192]*kernel[7]+tmp[193]*kernel[8];
				ans[93]<=tmp[92]*kernel[3]+tmp[93]*kernel[4]+tmp[94]*kernel[5]+tmp[192]*kernel[6]+tmp[193]*kernel[7]+tmp[194]*kernel[8];
				ans[94]<=tmp[93]*kernel[3]+tmp[94]*kernel[4]+tmp[95]*kernel[5]+tmp[193]*kernel[6]+tmp[194]*kernel[7]+tmp[195]*kernel[8];
				ans[95]<=tmp[94]*kernel[3]+tmp[95]*kernel[4]+tmp[96]*kernel[5]+tmp[194]*kernel[6]+tmp[195]*kernel[7]+tmp[196]*kernel[8];
				ans[96]<=tmp[95]*kernel[3]+tmp[96]*kernel[4]+tmp[97]*kernel[5]+tmp[195]*kernel[6]+tmp[196]*kernel[7]+tmp[197]*kernel[8];
				ans[97]<=tmp[96]*kernel[3]+tmp[97]*kernel[4]+tmp[98]*kernel[5]+tmp[196]*kernel[6]+tmp[197]*kernel[7]+tmp[198]*kernel[8];
				ans[98]<=tmp[97]*kernel[3]+tmp[98]*kernel[4]+tmp[99]*kernel[5]+tmp[197]*kernel[6]+tmp[198]*kernel[7]+tmp[199]*kernel[8];
				ans[99]<=tmp[98]*kernel[3]+tmp[99]*kernel[4]+tmp[198]*kernel[6]+tmp[199]*kernel[7];
				ans[100]<=tmp[0]*kernel[1]+tmp[1]*kernel[2]+tmp[100]*kernel[4]+tmp[101]*kernel[5]+tmp[200]*kernel[7]+tmp[201]*kernel[8];
				ans[101]<=tmp[0]*kernel[0]+tmp[1]*kernel[1]+tmp[2]*kernel[2]+tmp[100]*kernel[3]+tmp[101]*kernel[4]+tmp[102]*kernel[5]+tmp[200]*kernel[6]+tmp[201]*kernel[7]+tmp[202]*kernel[8];
				ans[102]<=tmp[1]*kernel[0]+tmp[2]*kernel[1]+tmp[3]*kernel[2]+tmp[101]*kernel[3]+tmp[102]*kernel[4]+tmp[103]*kernel[5]+tmp[201]*kernel[6]+tmp[202]*kernel[7]+tmp[203]*kernel[8];
				ans[103]<=tmp[2]*kernel[0]+tmp[3]*kernel[1]+tmp[4]*kernel[2]+tmp[102]*kernel[3]+tmp[103]*kernel[4]+tmp[104]*kernel[5]+tmp[202]*kernel[6]+tmp[203]*kernel[7]+tmp[204]*kernel[8];
				ans[104]<=tmp[3]*kernel[0]+tmp[4]*kernel[1]+tmp[5]*kernel[2]+tmp[103]*kernel[3]+tmp[104]*kernel[4]+tmp[105]*kernel[5]+tmp[203]*kernel[6]+tmp[204]*kernel[7]+tmp[205]*kernel[8];
				ans[105]<=tmp[4]*kernel[0]+tmp[5]*kernel[1]+tmp[6]*kernel[2]+tmp[104]*kernel[3]+tmp[105]*kernel[4]+tmp[106]*kernel[5]+tmp[204]*kernel[6]+tmp[205]*kernel[7]+tmp[206]*kernel[8];
				ans[106]<=tmp[5]*kernel[0]+tmp[6]*kernel[1]+tmp[7]*kernel[2]+tmp[105]*kernel[3]+tmp[106]*kernel[4]+tmp[107]*kernel[5]+tmp[205]*kernel[6]+tmp[206]*kernel[7]+tmp[207]*kernel[8];
				ans[107]<=tmp[6]*kernel[0]+tmp[7]*kernel[1]+tmp[8]*kernel[2]+tmp[106]*kernel[3]+tmp[107]*kernel[4]+tmp[108]*kernel[5]+tmp[206]*kernel[6]+tmp[207]*kernel[7]+tmp[208]*kernel[8];
				ans[108]<=tmp[7]*kernel[0]+tmp[8]*kernel[1]+tmp[9]*kernel[2]+tmp[107]*kernel[3]+tmp[108]*kernel[4]+tmp[109]*kernel[5]+tmp[207]*kernel[6]+tmp[208]*kernel[7]+tmp[209]*kernel[8];
				ans[109]<=tmp[8]*kernel[0]+tmp[9]*kernel[1]+tmp[10]*kernel[2]+tmp[108]*kernel[3]+tmp[109]*kernel[4]+tmp[110]*kernel[5]+tmp[208]*kernel[6]+tmp[209]*kernel[7]+tmp[210]*kernel[8];
				ans[110]<=tmp[9]*kernel[0]+tmp[10]*kernel[1]+tmp[11]*kernel[2]+tmp[109]*kernel[3]+tmp[110]*kernel[4]+tmp[111]*kernel[5]+tmp[209]*kernel[6]+tmp[210]*kernel[7]+tmp[211]*kernel[8];
				ans[111]<=tmp[10]*kernel[0]+tmp[11]*kernel[1]+tmp[12]*kernel[2]+tmp[110]*kernel[3]+tmp[111]*kernel[4]+tmp[112]*kernel[5]+tmp[210]*kernel[6]+tmp[211]*kernel[7]+tmp[212]*kernel[8];
				ans[112]<=tmp[11]*kernel[0]+tmp[12]*kernel[1]+tmp[13]*kernel[2]+tmp[111]*kernel[3]+tmp[112]*kernel[4]+tmp[113]*kernel[5]+tmp[211]*kernel[6]+tmp[212]*kernel[7]+tmp[213]*kernel[8];
				ans[113]<=tmp[12]*kernel[0]+tmp[13]*kernel[1]+tmp[14]*kernel[2]+tmp[112]*kernel[3]+tmp[113]*kernel[4]+tmp[114]*kernel[5]+tmp[212]*kernel[6]+tmp[213]*kernel[7]+tmp[214]*kernel[8];
				ans[114]<=tmp[13]*kernel[0]+tmp[14]*kernel[1]+tmp[15]*kernel[2]+tmp[113]*kernel[3]+tmp[114]*kernel[4]+tmp[115]*kernel[5]+tmp[213]*kernel[6]+tmp[214]*kernel[7]+tmp[215]*kernel[8];
				ans[115]<=tmp[14]*kernel[0]+tmp[15]*kernel[1]+tmp[16]*kernel[2]+tmp[114]*kernel[3]+tmp[115]*kernel[4]+tmp[116]*kernel[5]+tmp[214]*kernel[6]+tmp[215]*kernel[7]+tmp[216]*kernel[8];
				ans[116]<=tmp[15]*kernel[0]+tmp[16]*kernel[1]+tmp[17]*kernel[2]+tmp[115]*kernel[3]+tmp[116]*kernel[4]+tmp[117]*kernel[5]+tmp[215]*kernel[6]+tmp[216]*kernel[7]+tmp[217]*kernel[8];
				ans[117]<=tmp[16]*kernel[0]+tmp[17]*kernel[1]+tmp[18]*kernel[2]+tmp[116]*kernel[3]+tmp[117]*kernel[4]+tmp[118]*kernel[5]+tmp[216]*kernel[6]+tmp[217]*kernel[7]+tmp[218]*kernel[8];
				ans[118]<=tmp[17]*kernel[0]+tmp[18]*kernel[1]+tmp[19]*kernel[2]+tmp[117]*kernel[3]+tmp[118]*kernel[4]+tmp[119]*kernel[5]+tmp[217]*kernel[6]+tmp[218]*kernel[7]+tmp[219]*kernel[8];
				ans[119]<=tmp[18]*kernel[0]+tmp[19]*kernel[1]+tmp[20]*kernel[2]+tmp[118]*kernel[3]+tmp[119]*kernel[4]+tmp[120]*kernel[5]+tmp[218]*kernel[6]+tmp[219]*kernel[7]+tmp[220]*kernel[8];
				ans[120]<=tmp[19]*kernel[0]+tmp[20]*kernel[1]+tmp[21]*kernel[2]+tmp[119]*kernel[3]+tmp[120]*kernel[4]+tmp[121]*kernel[5]+tmp[219]*kernel[6]+tmp[220]*kernel[7]+tmp[221]*kernel[8];
				ans[121]<=tmp[20]*kernel[0]+tmp[21]*kernel[1]+tmp[22]*kernel[2]+tmp[120]*kernel[3]+tmp[121]*kernel[4]+tmp[122]*kernel[5]+tmp[220]*kernel[6]+tmp[221]*kernel[7]+tmp[222]*kernel[8];
				ans[122]<=tmp[21]*kernel[0]+tmp[22]*kernel[1]+tmp[23]*kernel[2]+tmp[121]*kernel[3]+tmp[122]*kernel[4]+tmp[123]*kernel[5]+tmp[221]*kernel[6]+tmp[222]*kernel[7]+tmp[223]*kernel[8];
				ans[123]<=tmp[22]*kernel[0]+tmp[23]*kernel[1]+tmp[24]*kernel[2]+tmp[122]*kernel[3]+tmp[123]*kernel[4]+tmp[124]*kernel[5]+tmp[222]*kernel[6]+tmp[223]*kernel[7]+tmp[224]*kernel[8];
				ans[124]<=tmp[23]*kernel[0]+tmp[24]*kernel[1]+tmp[25]*kernel[2]+tmp[123]*kernel[3]+tmp[124]*kernel[4]+tmp[125]*kernel[5]+tmp[223]*kernel[6]+tmp[224]*kernel[7]+tmp[225]*kernel[8];
				ans[125]<=tmp[24]*kernel[0]+tmp[25]*kernel[1]+tmp[26]*kernel[2]+tmp[124]*kernel[3]+tmp[125]*kernel[4]+tmp[126]*kernel[5]+tmp[224]*kernel[6]+tmp[225]*kernel[7]+tmp[226]*kernel[8];
				ans[126]<=tmp[25]*kernel[0]+tmp[26]*kernel[1]+tmp[27]*kernel[2]+tmp[125]*kernel[3]+tmp[126]*kernel[4]+tmp[127]*kernel[5]+tmp[225]*kernel[6]+tmp[226]*kernel[7]+tmp[227]*kernel[8];
				ans[127]<=tmp[26]*kernel[0]+tmp[27]*kernel[1]+tmp[28]*kernel[2]+tmp[126]*kernel[3]+tmp[127]*kernel[4]+tmp[128]*kernel[5]+tmp[226]*kernel[6]+tmp[227]*kernel[7]+tmp[228]*kernel[8];
				ans[128]<=tmp[27]*kernel[0]+tmp[28]*kernel[1]+tmp[29]*kernel[2]+tmp[127]*kernel[3]+tmp[128]*kernel[4]+tmp[129]*kernel[5]+tmp[227]*kernel[6]+tmp[228]*kernel[7]+tmp[229]*kernel[8];
				ans[129]<=tmp[28]*kernel[0]+tmp[29]*kernel[1]+tmp[30]*kernel[2]+tmp[128]*kernel[3]+tmp[129]*kernel[4]+tmp[130]*kernel[5]+tmp[228]*kernel[6]+tmp[229]*kernel[7]+tmp[230]*kernel[8];
				ans[130]<=tmp[29]*kernel[0]+tmp[30]*kernel[1]+tmp[31]*kernel[2]+tmp[129]*kernel[3]+tmp[130]*kernel[4]+tmp[131]*kernel[5]+tmp[229]*kernel[6]+tmp[230]*kernel[7]+tmp[231]*kernel[8];
				ans[131]<=tmp[30]*kernel[0]+tmp[31]*kernel[1]+tmp[32]*kernel[2]+tmp[130]*kernel[3]+tmp[131]*kernel[4]+tmp[132]*kernel[5]+tmp[230]*kernel[6]+tmp[231]*kernel[7]+tmp[232]*kernel[8];
				ans[132]<=tmp[31]*kernel[0]+tmp[32]*kernel[1]+tmp[33]*kernel[2]+tmp[131]*kernel[3]+tmp[132]*kernel[4]+tmp[133]*kernel[5]+tmp[231]*kernel[6]+tmp[232]*kernel[7]+tmp[233]*kernel[8];
				ans[133]<=tmp[32]*kernel[0]+tmp[33]*kernel[1]+tmp[34]*kernel[2]+tmp[132]*kernel[3]+tmp[133]*kernel[4]+tmp[134]*kernel[5]+tmp[232]*kernel[6]+tmp[233]*kernel[7]+tmp[234]*kernel[8];
				ans[134]<=tmp[33]*kernel[0]+tmp[34]*kernel[1]+tmp[35]*kernel[2]+tmp[133]*kernel[3]+tmp[134]*kernel[4]+tmp[135]*kernel[5]+tmp[233]*kernel[6]+tmp[234]*kernel[7]+tmp[235]*kernel[8];
				ans[135]<=tmp[34]*kernel[0]+tmp[35]*kernel[1]+tmp[36]*kernel[2]+tmp[134]*kernel[3]+tmp[135]*kernel[4]+tmp[136]*kernel[5]+tmp[234]*kernel[6]+tmp[235]*kernel[7]+tmp[236]*kernel[8];
				ans[136]<=tmp[35]*kernel[0]+tmp[36]*kernel[1]+tmp[37]*kernel[2]+tmp[135]*kernel[3]+tmp[136]*kernel[4]+tmp[137]*kernel[5]+tmp[235]*kernel[6]+tmp[236]*kernel[7]+tmp[237]*kernel[8];
				ans[137]<=tmp[36]*kernel[0]+tmp[37]*kernel[1]+tmp[38]*kernel[2]+tmp[136]*kernel[3]+tmp[137]*kernel[4]+tmp[138]*kernel[5]+tmp[236]*kernel[6]+tmp[237]*kernel[7]+tmp[238]*kernel[8];
				ans[138]<=tmp[37]*kernel[0]+tmp[38]*kernel[1]+tmp[39]*kernel[2]+tmp[137]*kernel[3]+tmp[138]*kernel[4]+tmp[139]*kernel[5]+tmp[237]*kernel[6]+tmp[238]*kernel[7]+tmp[239]*kernel[8];
				ans[139]<=tmp[38]*kernel[0]+tmp[39]*kernel[1]+tmp[40]*kernel[2]+tmp[138]*kernel[3]+tmp[139]*kernel[4]+tmp[140]*kernel[5]+tmp[238]*kernel[6]+tmp[239]*kernel[7]+tmp[240]*kernel[8];
				ans[140]<=tmp[39]*kernel[0]+tmp[40]*kernel[1]+tmp[41]*kernel[2]+tmp[139]*kernel[3]+tmp[140]*kernel[4]+tmp[141]*kernel[5]+tmp[239]*kernel[6]+tmp[240]*kernel[7]+tmp[241]*kernel[8];
				ans[141]<=tmp[40]*kernel[0]+tmp[41]*kernel[1]+tmp[42]*kernel[2]+tmp[140]*kernel[3]+tmp[141]*kernel[4]+tmp[142]*kernel[5]+tmp[240]*kernel[6]+tmp[241]*kernel[7]+tmp[242]*kernel[8];
				ans[142]<=tmp[41]*kernel[0]+tmp[42]*kernel[1]+tmp[43]*kernel[2]+tmp[141]*kernel[3]+tmp[142]*kernel[4]+tmp[143]*kernel[5]+tmp[241]*kernel[6]+tmp[242]*kernel[7]+tmp[243]*kernel[8];
				ans[143]<=tmp[42]*kernel[0]+tmp[43]*kernel[1]+tmp[44]*kernel[2]+tmp[142]*kernel[3]+tmp[143]*kernel[4]+tmp[144]*kernel[5]+tmp[242]*kernel[6]+tmp[243]*kernel[7]+tmp[244]*kernel[8];
				ans[144]<=tmp[43]*kernel[0]+tmp[44]*kernel[1]+tmp[45]*kernel[2]+tmp[143]*kernel[3]+tmp[144]*kernel[4]+tmp[145]*kernel[5]+tmp[243]*kernel[6]+tmp[244]*kernel[7]+tmp[245]*kernel[8];
				ans[145]<=tmp[44]*kernel[0]+tmp[45]*kernel[1]+tmp[46]*kernel[2]+tmp[144]*kernel[3]+tmp[145]*kernel[4]+tmp[146]*kernel[5]+tmp[244]*kernel[6]+tmp[245]*kernel[7]+tmp[246]*kernel[8];
				ans[146]<=tmp[45]*kernel[0]+tmp[46]*kernel[1]+tmp[47]*kernel[2]+tmp[145]*kernel[3]+tmp[146]*kernel[4]+tmp[147]*kernel[5]+tmp[245]*kernel[6]+tmp[246]*kernel[7]+tmp[247]*kernel[8];
				ans[147]<=tmp[46]*kernel[0]+tmp[47]*kernel[1]+tmp[48]*kernel[2]+tmp[146]*kernel[3]+tmp[147]*kernel[4]+tmp[148]*kernel[5]+tmp[246]*kernel[6]+tmp[247]*kernel[7]+tmp[248]*kernel[8];
				ans[148]<=tmp[47]*kernel[0]+tmp[48]*kernel[1]+tmp[49]*kernel[2]+tmp[147]*kernel[3]+tmp[148]*kernel[4]+tmp[149]*kernel[5]+tmp[247]*kernel[6]+tmp[248]*kernel[7]+tmp[249]*kernel[8];
				ans[149]<=tmp[48]*kernel[0]+tmp[49]*kernel[1]+tmp[50]*kernel[2]+tmp[148]*kernel[3]+tmp[149]*kernel[4]+tmp[150]*kernel[5]+tmp[248]*kernel[6]+tmp[249]*kernel[7]+tmp[250]*kernel[8];
				ans[150]<=tmp[49]*kernel[0]+tmp[50]*kernel[1]+tmp[51]*kernel[2]+tmp[149]*kernel[3]+tmp[150]*kernel[4]+tmp[151]*kernel[5]+tmp[249]*kernel[6]+tmp[250]*kernel[7]+tmp[251]*kernel[8];
				ans[151]<=tmp[50]*kernel[0]+tmp[51]*kernel[1]+tmp[52]*kernel[2]+tmp[150]*kernel[3]+tmp[151]*kernel[4]+tmp[152]*kernel[5]+tmp[250]*kernel[6]+tmp[251]*kernel[7]+tmp[252]*kernel[8];
				ans[152]<=tmp[51]*kernel[0]+tmp[52]*kernel[1]+tmp[53]*kernel[2]+tmp[151]*kernel[3]+tmp[152]*kernel[4]+tmp[153]*kernel[5]+tmp[251]*kernel[6]+tmp[252]*kernel[7]+tmp[253]*kernel[8];
				ans[153]<=tmp[52]*kernel[0]+tmp[53]*kernel[1]+tmp[54]*kernel[2]+tmp[152]*kernel[3]+tmp[153]*kernel[4]+tmp[154]*kernel[5]+tmp[252]*kernel[6]+tmp[253]*kernel[7]+tmp[254]*kernel[8];
				ans[154]<=tmp[53]*kernel[0]+tmp[54]*kernel[1]+tmp[55]*kernel[2]+tmp[153]*kernel[3]+tmp[154]*kernel[4]+tmp[155]*kernel[5]+tmp[253]*kernel[6]+tmp[254]*kernel[7]+tmp[255]*kernel[8];
				ans[155]<=tmp[54]*kernel[0]+tmp[55]*kernel[1]+tmp[56]*kernel[2]+tmp[154]*kernel[3]+tmp[155]*kernel[4]+tmp[156]*kernel[5]+tmp[254]*kernel[6]+tmp[255]*kernel[7]+tmp[256]*kernel[8];
				ans[156]<=tmp[55]*kernel[0]+tmp[56]*kernel[1]+tmp[57]*kernel[2]+tmp[155]*kernel[3]+tmp[156]*kernel[4]+tmp[157]*kernel[5]+tmp[255]*kernel[6]+tmp[256]*kernel[7]+tmp[257]*kernel[8];
				ans[157]<=tmp[56]*kernel[0]+tmp[57]*kernel[1]+tmp[58]*kernel[2]+tmp[156]*kernel[3]+tmp[157]*kernel[4]+tmp[158]*kernel[5]+tmp[256]*kernel[6]+tmp[257]*kernel[7]+tmp[258]*kernel[8];
				ans[158]<=tmp[57]*kernel[0]+tmp[58]*kernel[1]+tmp[59]*kernel[2]+tmp[157]*kernel[3]+tmp[158]*kernel[4]+tmp[159]*kernel[5]+tmp[257]*kernel[6]+tmp[258]*kernel[7]+tmp[259]*kernel[8];
				ans[159]<=tmp[58]*kernel[0]+tmp[59]*kernel[1]+tmp[60]*kernel[2]+tmp[158]*kernel[3]+tmp[159]*kernel[4]+tmp[160]*kernel[5]+tmp[258]*kernel[6]+tmp[259]*kernel[7]+tmp[260]*kernel[8];
				ans[160]<=tmp[59]*kernel[0]+tmp[60]*kernel[1]+tmp[61]*kernel[2]+tmp[159]*kernel[3]+tmp[160]*kernel[4]+tmp[161]*kernel[5]+tmp[259]*kernel[6]+tmp[260]*kernel[7]+tmp[261]*kernel[8];
				ans[161]<=tmp[60]*kernel[0]+tmp[61]*kernel[1]+tmp[62]*kernel[2]+tmp[160]*kernel[3]+tmp[161]*kernel[4]+tmp[162]*kernel[5]+tmp[260]*kernel[6]+tmp[261]*kernel[7]+tmp[262]*kernel[8];
				ans[162]<=tmp[61]*kernel[0]+tmp[62]*kernel[1]+tmp[63]*kernel[2]+tmp[161]*kernel[3]+tmp[162]*kernel[4]+tmp[163]*kernel[5]+tmp[261]*kernel[6]+tmp[262]*kernel[7]+tmp[263]*kernel[8];
				ans[163]<=tmp[62]*kernel[0]+tmp[63]*kernel[1]+tmp[64]*kernel[2]+tmp[162]*kernel[3]+tmp[163]*kernel[4]+tmp[164]*kernel[5]+tmp[262]*kernel[6]+tmp[263]*kernel[7]+tmp[264]*kernel[8];
				ans[164]<=tmp[63]*kernel[0]+tmp[64]*kernel[1]+tmp[65]*kernel[2]+tmp[163]*kernel[3]+tmp[164]*kernel[4]+tmp[165]*kernel[5]+tmp[263]*kernel[6]+tmp[264]*kernel[7]+tmp[265]*kernel[8];
				ans[165]<=tmp[64]*kernel[0]+tmp[65]*kernel[1]+tmp[66]*kernel[2]+tmp[164]*kernel[3]+tmp[165]*kernel[4]+tmp[166]*kernel[5]+tmp[264]*kernel[6]+tmp[265]*kernel[7]+tmp[266]*kernel[8];
				ans[166]<=tmp[65]*kernel[0]+tmp[66]*kernel[1]+tmp[67]*kernel[2]+tmp[165]*kernel[3]+tmp[166]*kernel[4]+tmp[167]*kernel[5]+tmp[265]*kernel[6]+tmp[266]*kernel[7]+tmp[267]*kernel[8];
				ans[167]<=tmp[66]*kernel[0]+tmp[67]*kernel[1]+tmp[68]*kernel[2]+tmp[166]*kernel[3]+tmp[167]*kernel[4]+tmp[168]*kernel[5]+tmp[266]*kernel[6]+tmp[267]*kernel[7]+tmp[268]*kernel[8];
				ans[168]<=tmp[67]*kernel[0]+tmp[68]*kernel[1]+tmp[69]*kernel[2]+tmp[167]*kernel[3]+tmp[168]*kernel[4]+tmp[169]*kernel[5]+tmp[267]*kernel[6]+tmp[268]*kernel[7]+tmp[269]*kernel[8];
				ans[169]<=tmp[68]*kernel[0]+tmp[69]*kernel[1]+tmp[70]*kernel[2]+tmp[168]*kernel[3]+tmp[169]*kernel[4]+tmp[170]*kernel[5]+tmp[268]*kernel[6]+tmp[269]*kernel[7]+tmp[270]*kernel[8];
				ans[170]<=tmp[69]*kernel[0]+tmp[70]*kernel[1]+tmp[71]*kernel[2]+tmp[169]*kernel[3]+tmp[170]*kernel[4]+tmp[171]*kernel[5]+tmp[269]*kernel[6]+tmp[270]*kernel[7]+tmp[271]*kernel[8];
				ans[171]<=tmp[70]*kernel[0]+tmp[71]*kernel[1]+tmp[72]*kernel[2]+tmp[170]*kernel[3]+tmp[171]*kernel[4]+tmp[172]*kernel[5]+tmp[270]*kernel[6]+tmp[271]*kernel[7]+tmp[272]*kernel[8];
				ans[172]<=tmp[71]*kernel[0]+tmp[72]*kernel[1]+tmp[73]*kernel[2]+tmp[171]*kernel[3]+tmp[172]*kernel[4]+tmp[173]*kernel[5]+tmp[271]*kernel[6]+tmp[272]*kernel[7]+tmp[273]*kernel[8];
				ans[173]<=tmp[72]*kernel[0]+tmp[73]*kernel[1]+tmp[74]*kernel[2]+tmp[172]*kernel[3]+tmp[173]*kernel[4]+tmp[174]*kernel[5]+tmp[272]*kernel[6]+tmp[273]*kernel[7]+tmp[274]*kernel[8];
				ans[174]<=tmp[73]*kernel[0]+tmp[74]*kernel[1]+tmp[75]*kernel[2]+tmp[173]*kernel[3]+tmp[174]*kernel[4]+tmp[175]*kernel[5]+tmp[273]*kernel[6]+tmp[274]*kernel[7]+tmp[275]*kernel[8];
				ans[175]<=tmp[74]*kernel[0]+tmp[75]*kernel[1]+tmp[76]*kernel[2]+tmp[174]*kernel[3]+tmp[175]*kernel[4]+tmp[176]*kernel[5]+tmp[274]*kernel[6]+tmp[275]*kernel[7]+tmp[276]*kernel[8];
				ans[176]<=tmp[75]*kernel[0]+tmp[76]*kernel[1]+tmp[77]*kernel[2]+tmp[175]*kernel[3]+tmp[176]*kernel[4]+tmp[177]*kernel[5]+tmp[275]*kernel[6]+tmp[276]*kernel[7]+tmp[277]*kernel[8];
				ans[177]<=tmp[76]*kernel[0]+tmp[77]*kernel[1]+tmp[78]*kernel[2]+tmp[176]*kernel[3]+tmp[177]*kernel[4]+tmp[178]*kernel[5]+tmp[276]*kernel[6]+tmp[277]*kernel[7]+tmp[278]*kernel[8];
				ans[178]<=tmp[77]*kernel[0]+tmp[78]*kernel[1]+tmp[79]*kernel[2]+tmp[177]*kernel[3]+tmp[178]*kernel[4]+tmp[179]*kernel[5]+tmp[277]*kernel[6]+tmp[278]*kernel[7]+tmp[279]*kernel[8];
				ans[179]<=tmp[78]*kernel[0]+tmp[79]*kernel[1]+tmp[80]*kernel[2]+tmp[178]*kernel[3]+tmp[179]*kernel[4]+tmp[180]*kernel[5]+tmp[278]*kernel[6]+tmp[279]*kernel[7]+tmp[280]*kernel[8];
				ans[180]<=tmp[79]*kernel[0]+tmp[80]*kernel[1]+tmp[81]*kernel[2]+tmp[179]*kernel[3]+tmp[180]*kernel[4]+tmp[181]*kernel[5]+tmp[279]*kernel[6]+tmp[280]*kernel[7]+tmp[281]*kernel[8];
				ans[181]<=tmp[80]*kernel[0]+tmp[81]*kernel[1]+tmp[82]*kernel[2]+tmp[180]*kernel[3]+tmp[181]*kernel[4]+tmp[182]*kernel[5]+tmp[280]*kernel[6]+tmp[281]*kernel[7]+tmp[282]*kernel[8];
				ans[182]<=tmp[81]*kernel[0]+tmp[82]*kernel[1]+tmp[83]*kernel[2]+tmp[181]*kernel[3]+tmp[182]*kernel[4]+tmp[183]*kernel[5]+tmp[281]*kernel[6]+tmp[282]*kernel[7]+tmp[283]*kernel[8];
				ans[183]<=tmp[82]*kernel[0]+tmp[83]*kernel[1]+tmp[84]*kernel[2]+tmp[182]*kernel[3]+tmp[183]*kernel[4]+tmp[184]*kernel[5]+tmp[282]*kernel[6]+tmp[283]*kernel[7]+tmp[284]*kernel[8];
				ans[184]<=tmp[83]*kernel[0]+tmp[84]*kernel[1]+tmp[85]*kernel[2]+tmp[183]*kernel[3]+tmp[184]*kernel[4]+tmp[185]*kernel[5]+tmp[283]*kernel[6]+tmp[284]*kernel[7]+tmp[285]*kernel[8];
				ans[185]<=tmp[84]*kernel[0]+tmp[85]*kernel[1]+tmp[86]*kernel[2]+tmp[184]*kernel[3]+tmp[185]*kernel[4]+tmp[186]*kernel[5]+tmp[284]*kernel[6]+tmp[285]*kernel[7]+tmp[286]*kernel[8];
				ans[186]<=tmp[85]*kernel[0]+tmp[86]*kernel[1]+tmp[87]*kernel[2]+tmp[185]*kernel[3]+tmp[186]*kernel[4]+tmp[187]*kernel[5]+tmp[285]*kernel[6]+tmp[286]*kernel[7]+tmp[287]*kernel[8];
				ans[187]<=tmp[86]*kernel[0]+tmp[87]*kernel[1]+tmp[88]*kernel[2]+tmp[186]*kernel[3]+tmp[187]*kernel[4]+tmp[188]*kernel[5]+tmp[286]*kernel[6]+tmp[287]*kernel[7]+tmp[288]*kernel[8];
				ans[188]<=tmp[87]*kernel[0]+tmp[88]*kernel[1]+tmp[89]*kernel[2]+tmp[187]*kernel[3]+tmp[188]*kernel[4]+tmp[189]*kernel[5]+tmp[287]*kernel[6]+tmp[288]*kernel[7]+tmp[289]*kernel[8];
				ans[189]<=tmp[88]*kernel[0]+tmp[89]*kernel[1]+tmp[90]*kernel[2]+tmp[188]*kernel[3]+tmp[189]*kernel[4]+tmp[190]*kernel[5]+tmp[288]*kernel[6]+tmp[289]*kernel[7]+tmp[290]*kernel[8];
				ans[190]<=tmp[89]*kernel[0]+tmp[90]*kernel[1]+tmp[91]*kernel[2]+tmp[189]*kernel[3]+tmp[190]*kernel[4]+tmp[191]*kernel[5]+tmp[289]*kernel[6]+tmp[290]*kernel[7]+tmp[291]*kernel[8];
				ans[191]<=tmp[90]*kernel[0]+tmp[91]*kernel[1]+tmp[92]*kernel[2]+tmp[190]*kernel[3]+tmp[191]*kernel[4]+tmp[192]*kernel[5]+tmp[290]*kernel[6]+tmp[291]*kernel[7]+tmp[292]*kernel[8];
				ans[192]<=tmp[91]*kernel[0]+tmp[92]*kernel[1]+tmp[93]*kernel[2]+tmp[191]*kernel[3]+tmp[192]*kernel[4]+tmp[193]*kernel[5]+tmp[291]*kernel[6]+tmp[292]*kernel[7]+tmp[293]*kernel[8];
				ans[193]<=tmp[92]*kernel[0]+tmp[93]*kernel[1]+tmp[94]*kernel[2]+tmp[192]*kernel[3]+tmp[193]*kernel[4]+tmp[194]*kernel[5]+tmp[292]*kernel[6]+tmp[293]*kernel[7]+tmp[294]*kernel[8];
				ans[194]<=tmp[93]*kernel[0]+tmp[94]*kernel[1]+tmp[95]*kernel[2]+tmp[193]*kernel[3]+tmp[194]*kernel[4]+tmp[195]*kernel[5]+tmp[293]*kernel[6]+tmp[294]*kernel[7]+tmp[295]*kernel[8];
				ans[195]<=tmp[94]*kernel[0]+tmp[95]*kernel[1]+tmp[96]*kernel[2]+tmp[194]*kernel[3]+tmp[195]*kernel[4]+tmp[196]*kernel[5]+tmp[294]*kernel[6]+tmp[295]*kernel[7]+tmp[296]*kernel[8];
				ans[196]<=tmp[95]*kernel[0]+tmp[96]*kernel[1]+tmp[97]*kernel[2]+tmp[195]*kernel[3]+tmp[196]*kernel[4]+tmp[197]*kernel[5]+tmp[295]*kernel[6]+tmp[296]*kernel[7]+tmp[297]*kernel[8];
				ans[197]<=tmp[96]*kernel[0]+tmp[97]*kernel[1]+tmp[98]*kernel[2]+tmp[196]*kernel[3]+tmp[197]*kernel[4]+tmp[198]*kernel[5]+tmp[296]*kernel[6]+tmp[297]*kernel[7]+tmp[298]*kernel[8];
				ans[198]<=tmp[97]*kernel[0]+tmp[98]*kernel[1]+tmp[99]*kernel[2]+tmp[197]*kernel[3]+tmp[198]*kernel[4]+tmp[199]*kernel[5]+tmp[297]*kernel[6]+tmp[298]*kernel[7]+tmp[299]*kernel[8];
				ans[199]<=tmp[98]*kernel[0]+tmp[99]*kernel[1]+tmp[198]*kernel[3]+tmp[199]*kernel[4]+tmp[298]*kernel[6]+tmp[299]*kernel[7];
				ans[200]<=tmp[100]*kernel[1]+tmp[101]*kernel[2]+tmp[200]*kernel[4]+tmp[201]*kernel[5]+tmp[300]*kernel[7]+tmp[301]*kernel[8];
				ans[201]<=tmp[100]*kernel[0]+tmp[101]*kernel[1]+tmp[102]*kernel[2]+tmp[200]*kernel[3]+tmp[201]*kernel[4]+tmp[202]*kernel[5]+tmp[300]*kernel[6]+tmp[301]*kernel[7]+tmp[302]*kernel[8];
				ans[202]<=tmp[101]*kernel[0]+tmp[102]*kernel[1]+tmp[103]*kernel[2]+tmp[201]*kernel[3]+tmp[202]*kernel[4]+tmp[203]*kernel[5]+tmp[301]*kernel[6]+tmp[302]*kernel[7]+tmp[303]*kernel[8];
				ans[203]<=tmp[102]*kernel[0]+tmp[103]*kernel[1]+tmp[104]*kernel[2]+tmp[202]*kernel[3]+tmp[203]*kernel[4]+tmp[204]*kernel[5]+tmp[302]*kernel[6]+tmp[303]*kernel[7]+tmp[304]*kernel[8];
				ans[204]<=tmp[103]*kernel[0]+tmp[104]*kernel[1]+tmp[105]*kernel[2]+tmp[203]*kernel[3]+tmp[204]*kernel[4]+tmp[205]*kernel[5]+tmp[303]*kernel[6]+tmp[304]*kernel[7]+tmp[305]*kernel[8];
				ans[205]<=tmp[104]*kernel[0]+tmp[105]*kernel[1]+tmp[106]*kernel[2]+tmp[204]*kernel[3]+tmp[205]*kernel[4]+tmp[206]*kernel[5]+tmp[304]*kernel[6]+tmp[305]*kernel[7]+tmp[306]*kernel[8];
				ans[206]<=tmp[105]*kernel[0]+tmp[106]*kernel[1]+tmp[107]*kernel[2]+tmp[205]*kernel[3]+tmp[206]*kernel[4]+tmp[207]*kernel[5]+tmp[305]*kernel[6]+tmp[306]*kernel[7]+tmp[307]*kernel[8];
				ans[207]<=tmp[106]*kernel[0]+tmp[107]*kernel[1]+tmp[108]*kernel[2]+tmp[206]*kernel[3]+tmp[207]*kernel[4]+tmp[208]*kernel[5]+tmp[306]*kernel[6]+tmp[307]*kernel[7]+tmp[308]*kernel[8];
				ans[208]<=tmp[107]*kernel[0]+tmp[108]*kernel[1]+tmp[109]*kernel[2]+tmp[207]*kernel[3]+tmp[208]*kernel[4]+tmp[209]*kernel[5]+tmp[307]*kernel[6]+tmp[308]*kernel[7]+tmp[309]*kernel[8];
				ans[209]<=tmp[108]*kernel[0]+tmp[109]*kernel[1]+tmp[110]*kernel[2]+tmp[208]*kernel[3]+tmp[209]*kernel[4]+tmp[210]*kernel[5]+tmp[308]*kernel[6]+tmp[309]*kernel[7]+tmp[310]*kernel[8];
				ans[210]<=tmp[109]*kernel[0]+tmp[110]*kernel[1]+tmp[111]*kernel[2]+tmp[209]*kernel[3]+tmp[210]*kernel[4]+tmp[211]*kernel[5]+tmp[309]*kernel[6]+tmp[310]*kernel[7]+tmp[311]*kernel[8];
				ans[211]<=tmp[110]*kernel[0]+tmp[111]*kernel[1]+tmp[112]*kernel[2]+tmp[210]*kernel[3]+tmp[211]*kernel[4]+tmp[212]*kernel[5]+tmp[310]*kernel[6]+tmp[311]*kernel[7]+tmp[312]*kernel[8];
				ans[212]<=tmp[111]*kernel[0]+tmp[112]*kernel[1]+tmp[113]*kernel[2]+tmp[211]*kernel[3]+tmp[212]*kernel[4]+tmp[213]*kernel[5]+tmp[311]*kernel[6]+tmp[312]*kernel[7]+tmp[313]*kernel[8];
				ans[213]<=tmp[112]*kernel[0]+tmp[113]*kernel[1]+tmp[114]*kernel[2]+tmp[212]*kernel[3]+tmp[213]*kernel[4]+tmp[214]*kernel[5]+tmp[312]*kernel[6]+tmp[313]*kernel[7]+tmp[314]*kernel[8];
				ans[214]<=tmp[113]*kernel[0]+tmp[114]*kernel[1]+tmp[115]*kernel[2]+tmp[213]*kernel[3]+tmp[214]*kernel[4]+tmp[215]*kernel[5]+tmp[313]*kernel[6]+tmp[314]*kernel[7]+tmp[315]*kernel[8];
				ans[215]<=tmp[114]*kernel[0]+tmp[115]*kernel[1]+tmp[116]*kernel[2]+tmp[214]*kernel[3]+tmp[215]*kernel[4]+tmp[216]*kernel[5]+tmp[314]*kernel[6]+tmp[315]*kernel[7]+tmp[316]*kernel[8];
				ans[216]<=tmp[115]*kernel[0]+tmp[116]*kernel[1]+tmp[117]*kernel[2]+tmp[215]*kernel[3]+tmp[216]*kernel[4]+tmp[217]*kernel[5]+tmp[315]*kernel[6]+tmp[316]*kernel[7]+tmp[317]*kernel[8];
				ans[217]<=tmp[116]*kernel[0]+tmp[117]*kernel[1]+tmp[118]*kernel[2]+tmp[216]*kernel[3]+tmp[217]*kernel[4]+tmp[218]*kernel[5]+tmp[316]*kernel[6]+tmp[317]*kernel[7]+tmp[318]*kernel[8];
				ans[218]<=tmp[117]*kernel[0]+tmp[118]*kernel[1]+tmp[119]*kernel[2]+tmp[217]*kernel[3]+tmp[218]*kernel[4]+tmp[219]*kernel[5]+tmp[317]*kernel[6]+tmp[318]*kernel[7]+tmp[319]*kernel[8];
				ans[219]<=tmp[118]*kernel[0]+tmp[119]*kernel[1]+tmp[120]*kernel[2]+tmp[218]*kernel[3]+tmp[219]*kernel[4]+tmp[220]*kernel[5]+tmp[318]*kernel[6]+tmp[319]*kernel[7]+tmp[320]*kernel[8];
				ans[220]<=tmp[119]*kernel[0]+tmp[120]*kernel[1]+tmp[121]*kernel[2]+tmp[219]*kernel[3]+tmp[220]*kernel[4]+tmp[221]*kernel[5]+tmp[319]*kernel[6]+tmp[320]*kernel[7]+tmp[321]*kernel[8];
				ans[221]<=tmp[120]*kernel[0]+tmp[121]*kernel[1]+tmp[122]*kernel[2]+tmp[220]*kernel[3]+tmp[221]*kernel[4]+tmp[222]*kernel[5]+tmp[320]*kernel[6]+tmp[321]*kernel[7]+tmp[322]*kernel[8];
				ans[222]<=tmp[121]*kernel[0]+tmp[122]*kernel[1]+tmp[123]*kernel[2]+tmp[221]*kernel[3]+tmp[222]*kernel[4]+tmp[223]*kernel[5]+tmp[321]*kernel[6]+tmp[322]*kernel[7]+tmp[323]*kernel[8];
				ans[223]<=tmp[122]*kernel[0]+tmp[123]*kernel[1]+tmp[124]*kernel[2]+tmp[222]*kernel[3]+tmp[223]*kernel[4]+tmp[224]*kernel[5]+tmp[322]*kernel[6]+tmp[323]*kernel[7]+tmp[324]*kernel[8];
				ans[224]<=tmp[123]*kernel[0]+tmp[124]*kernel[1]+tmp[125]*kernel[2]+tmp[223]*kernel[3]+tmp[224]*kernel[4]+tmp[225]*kernel[5]+tmp[323]*kernel[6]+tmp[324]*kernel[7]+tmp[325]*kernel[8];
				ans[225]<=tmp[124]*kernel[0]+tmp[125]*kernel[1]+tmp[126]*kernel[2]+tmp[224]*kernel[3]+tmp[225]*kernel[4]+tmp[226]*kernel[5]+tmp[324]*kernel[6]+tmp[325]*kernel[7]+tmp[326]*kernel[8];
				ans[226]<=tmp[125]*kernel[0]+tmp[126]*kernel[1]+tmp[127]*kernel[2]+tmp[225]*kernel[3]+tmp[226]*kernel[4]+tmp[227]*kernel[5]+tmp[325]*kernel[6]+tmp[326]*kernel[7]+tmp[327]*kernel[8];
				ans[227]<=tmp[126]*kernel[0]+tmp[127]*kernel[1]+tmp[128]*kernel[2]+tmp[226]*kernel[3]+tmp[227]*kernel[4]+tmp[228]*kernel[5]+tmp[326]*kernel[6]+tmp[327]*kernel[7]+tmp[328]*kernel[8];
				ans[228]<=tmp[127]*kernel[0]+tmp[128]*kernel[1]+tmp[129]*kernel[2]+tmp[227]*kernel[3]+tmp[228]*kernel[4]+tmp[229]*kernel[5]+tmp[327]*kernel[6]+tmp[328]*kernel[7]+tmp[329]*kernel[8];
				ans[229]<=tmp[128]*kernel[0]+tmp[129]*kernel[1]+tmp[130]*kernel[2]+tmp[228]*kernel[3]+tmp[229]*kernel[4]+tmp[230]*kernel[5]+tmp[328]*kernel[6]+tmp[329]*kernel[7]+tmp[330]*kernel[8];
				ans[230]<=tmp[129]*kernel[0]+tmp[130]*kernel[1]+tmp[131]*kernel[2]+tmp[229]*kernel[3]+tmp[230]*kernel[4]+tmp[231]*kernel[5]+tmp[329]*kernel[6]+tmp[330]*kernel[7]+tmp[331]*kernel[8];
				ans[231]<=tmp[130]*kernel[0]+tmp[131]*kernel[1]+tmp[132]*kernel[2]+tmp[230]*kernel[3]+tmp[231]*kernel[4]+tmp[232]*kernel[5]+tmp[330]*kernel[6]+tmp[331]*kernel[7]+tmp[332]*kernel[8];
				ans[232]<=tmp[131]*kernel[0]+tmp[132]*kernel[1]+tmp[133]*kernel[2]+tmp[231]*kernel[3]+tmp[232]*kernel[4]+tmp[233]*kernel[5]+tmp[331]*kernel[6]+tmp[332]*kernel[7]+tmp[333]*kernel[8];
				ans[233]<=tmp[132]*kernel[0]+tmp[133]*kernel[1]+tmp[134]*kernel[2]+tmp[232]*kernel[3]+tmp[233]*kernel[4]+tmp[234]*kernel[5]+tmp[332]*kernel[6]+tmp[333]*kernel[7]+tmp[334]*kernel[8];
				ans[234]<=tmp[133]*kernel[0]+tmp[134]*kernel[1]+tmp[135]*kernel[2]+tmp[233]*kernel[3]+tmp[234]*kernel[4]+tmp[235]*kernel[5]+tmp[333]*kernel[6]+tmp[334]*kernel[7]+tmp[335]*kernel[8];
				ans[235]<=tmp[134]*kernel[0]+tmp[135]*kernel[1]+tmp[136]*kernel[2]+tmp[234]*kernel[3]+tmp[235]*kernel[4]+tmp[236]*kernel[5]+tmp[334]*kernel[6]+tmp[335]*kernel[7]+tmp[336]*kernel[8];
				ans[236]<=tmp[135]*kernel[0]+tmp[136]*kernel[1]+tmp[137]*kernel[2]+tmp[235]*kernel[3]+tmp[236]*kernel[4]+tmp[237]*kernel[5]+tmp[335]*kernel[6]+tmp[336]*kernel[7]+tmp[337]*kernel[8];
				ans[237]<=tmp[136]*kernel[0]+tmp[137]*kernel[1]+tmp[138]*kernel[2]+tmp[236]*kernel[3]+tmp[237]*kernel[4]+tmp[238]*kernel[5]+tmp[336]*kernel[6]+tmp[337]*kernel[7]+tmp[338]*kernel[8];
				ans[238]<=tmp[137]*kernel[0]+tmp[138]*kernel[1]+tmp[139]*kernel[2]+tmp[237]*kernel[3]+tmp[238]*kernel[4]+tmp[239]*kernel[5]+tmp[337]*kernel[6]+tmp[338]*kernel[7]+tmp[339]*kernel[8];
				ans[239]<=tmp[138]*kernel[0]+tmp[139]*kernel[1]+tmp[140]*kernel[2]+tmp[238]*kernel[3]+tmp[239]*kernel[4]+tmp[240]*kernel[5]+tmp[338]*kernel[6]+tmp[339]*kernel[7]+tmp[340]*kernel[8];
				ans[240]<=tmp[139]*kernel[0]+tmp[140]*kernel[1]+tmp[141]*kernel[2]+tmp[239]*kernel[3]+tmp[240]*kernel[4]+tmp[241]*kernel[5]+tmp[339]*kernel[6]+tmp[340]*kernel[7]+tmp[341]*kernel[8];
				ans[241]<=tmp[140]*kernel[0]+tmp[141]*kernel[1]+tmp[142]*kernel[2]+tmp[240]*kernel[3]+tmp[241]*kernel[4]+tmp[242]*kernel[5]+tmp[340]*kernel[6]+tmp[341]*kernel[7]+tmp[342]*kernel[8];
				ans[242]<=tmp[141]*kernel[0]+tmp[142]*kernel[1]+tmp[143]*kernel[2]+tmp[241]*kernel[3]+tmp[242]*kernel[4]+tmp[243]*kernel[5]+tmp[341]*kernel[6]+tmp[342]*kernel[7]+tmp[343]*kernel[8];
				ans[243]<=tmp[142]*kernel[0]+tmp[143]*kernel[1]+tmp[144]*kernel[2]+tmp[242]*kernel[3]+tmp[243]*kernel[4]+tmp[244]*kernel[5]+tmp[342]*kernel[6]+tmp[343]*kernel[7]+tmp[344]*kernel[8];
				ans[244]<=tmp[143]*kernel[0]+tmp[144]*kernel[1]+tmp[145]*kernel[2]+tmp[243]*kernel[3]+tmp[244]*kernel[4]+tmp[245]*kernel[5]+tmp[343]*kernel[6]+tmp[344]*kernel[7]+tmp[345]*kernel[8];
				ans[245]<=tmp[144]*kernel[0]+tmp[145]*kernel[1]+tmp[146]*kernel[2]+tmp[244]*kernel[3]+tmp[245]*kernel[4]+tmp[246]*kernel[5]+tmp[344]*kernel[6]+tmp[345]*kernel[7]+tmp[346]*kernel[8];
				ans[246]<=tmp[145]*kernel[0]+tmp[146]*kernel[1]+tmp[147]*kernel[2]+tmp[245]*kernel[3]+tmp[246]*kernel[4]+tmp[247]*kernel[5]+tmp[345]*kernel[6]+tmp[346]*kernel[7]+tmp[347]*kernel[8];
				ans[247]<=tmp[146]*kernel[0]+tmp[147]*kernel[1]+tmp[148]*kernel[2]+tmp[246]*kernel[3]+tmp[247]*kernel[4]+tmp[248]*kernel[5]+tmp[346]*kernel[6]+tmp[347]*kernel[7]+tmp[348]*kernel[8];
				ans[248]<=tmp[147]*kernel[0]+tmp[148]*kernel[1]+tmp[149]*kernel[2]+tmp[247]*kernel[3]+tmp[248]*kernel[4]+tmp[249]*kernel[5]+tmp[347]*kernel[6]+tmp[348]*kernel[7]+tmp[349]*kernel[8];
				ans[249]<=tmp[148]*kernel[0]+tmp[149]*kernel[1]+tmp[150]*kernel[2]+tmp[248]*kernel[3]+tmp[249]*kernel[4]+tmp[250]*kernel[5]+tmp[348]*kernel[6]+tmp[349]*kernel[7]+tmp[350]*kernel[8];
				ans[250]<=tmp[149]*kernel[0]+tmp[150]*kernel[1]+tmp[151]*kernel[2]+tmp[249]*kernel[3]+tmp[250]*kernel[4]+tmp[251]*kernel[5]+tmp[349]*kernel[6]+tmp[350]*kernel[7]+tmp[351]*kernel[8];
				ans[251]<=tmp[150]*kernel[0]+tmp[151]*kernel[1]+tmp[152]*kernel[2]+tmp[250]*kernel[3]+tmp[251]*kernel[4]+tmp[252]*kernel[5]+tmp[350]*kernel[6]+tmp[351]*kernel[7]+tmp[352]*kernel[8];
				ans[252]<=tmp[151]*kernel[0]+tmp[152]*kernel[1]+tmp[153]*kernel[2]+tmp[251]*kernel[3]+tmp[252]*kernel[4]+tmp[253]*kernel[5]+tmp[351]*kernel[6]+tmp[352]*kernel[7]+tmp[353]*kernel[8];
				ans[253]<=tmp[152]*kernel[0]+tmp[153]*kernel[1]+tmp[154]*kernel[2]+tmp[252]*kernel[3]+tmp[253]*kernel[4]+tmp[254]*kernel[5]+tmp[352]*kernel[6]+tmp[353]*kernel[7]+tmp[354]*kernel[8];
				ans[254]<=tmp[153]*kernel[0]+tmp[154]*kernel[1]+tmp[155]*kernel[2]+tmp[253]*kernel[3]+tmp[254]*kernel[4]+tmp[255]*kernel[5]+tmp[353]*kernel[6]+tmp[354]*kernel[7]+tmp[355]*kernel[8];
				ans[255]<=tmp[154]*kernel[0]+tmp[155]*kernel[1]+tmp[156]*kernel[2]+tmp[254]*kernel[3]+tmp[255]*kernel[4]+tmp[256]*kernel[5]+tmp[354]*kernel[6]+tmp[355]*kernel[7]+tmp[356]*kernel[8];
				ans[256]<=tmp[155]*kernel[0]+tmp[156]*kernel[1]+tmp[157]*kernel[2]+tmp[255]*kernel[3]+tmp[256]*kernel[4]+tmp[257]*kernel[5]+tmp[355]*kernel[6]+tmp[356]*kernel[7]+tmp[357]*kernel[8];
				ans[257]<=tmp[156]*kernel[0]+tmp[157]*kernel[1]+tmp[158]*kernel[2]+tmp[256]*kernel[3]+tmp[257]*kernel[4]+tmp[258]*kernel[5]+tmp[356]*kernel[6]+tmp[357]*kernel[7]+tmp[358]*kernel[8];
				ans[258]<=tmp[157]*kernel[0]+tmp[158]*kernel[1]+tmp[159]*kernel[2]+tmp[257]*kernel[3]+tmp[258]*kernel[4]+tmp[259]*kernel[5]+tmp[357]*kernel[6]+tmp[358]*kernel[7]+tmp[359]*kernel[8];
				ans[259]<=tmp[158]*kernel[0]+tmp[159]*kernel[1]+tmp[160]*kernel[2]+tmp[258]*kernel[3]+tmp[259]*kernel[4]+tmp[260]*kernel[5]+tmp[358]*kernel[6]+tmp[359]*kernel[7]+tmp[360]*kernel[8];
				ans[260]<=tmp[159]*kernel[0]+tmp[160]*kernel[1]+tmp[161]*kernel[2]+tmp[259]*kernel[3]+tmp[260]*kernel[4]+tmp[261]*kernel[5]+tmp[359]*kernel[6]+tmp[360]*kernel[7]+tmp[361]*kernel[8];
				ans[261]<=tmp[160]*kernel[0]+tmp[161]*kernel[1]+tmp[162]*kernel[2]+tmp[260]*kernel[3]+tmp[261]*kernel[4]+tmp[262]*kernel[5]+tmp[360]*kernel[6]+tmp[361]*kernel[7]+tmp[362]*kernel[8];
				ans[262]<=tmp[161]*kernel[0]+tmp[162]*kernel[1]+tmp[163]*kernel[2]+tmp[261]*kernel[3]+tmp[262]*kernel[4]+tmp[263]*kernel[5]+tmp[361]*kernel[6]+tmp[362]*kernel[7]+tmp[363]*kernel[8];
				ans[263]<=tmp[162]*kernel[0]+tmp[163]*kernel[1]+tmp[164]*kernel[2]+tmp[262]*kernel[3]+tmp[263]*kernel[4]+tmp[264]*kernel[5]+tmp[362]*kernel[6]+tmp[363]*kernel[7]+tmp[364]*kernel[8];
				ans[264]<=tmp[163]*kernel[0]+tmp[164]*kernel[1]+tmp[165]*kernel[2]+tmp[263]*kernel[3]+tmp[264]*kernel[4]+tmp[265]*kernel[5]+tmp[363]*kernel[6]+tmp[364]*kernel[7]+tmp[365]*kernel[8];
				ans[265]<=tmp[164]*kernel[0]+tmp[165]*kernel[1]+tmp[166]*kernel[2]+tmp[264]*kernel[3]+tmp[265]*kernel[4]+tmp[266]*kernel[5]+tmp[364]*kernel[6]+tmp[365]*kernel[7]+tmp[366]*kernel[8];
				ans[266]<=tmp[165]*kernel[0]+tmp[166]*kernel[1]+tmp[167]*kernel[2]+tmp[265]*kernel[3]+tmp[266]*kernel[4]+tmp[267]*kernel[5]+tmp[365]*kernel[6]+tmp[366]*kernel[7]+tmp[367]*kernel[8];
				ans[267]<=tmp[166]*kernel[0]+tmp[167]*kernel[1]+tmp[168]*kernel[2]+tmp[266]*kernel[3]+tmp[267]*kernel[4]+tmp[268]*kernel[5]+tmp[366]*kernel[6]+tmp[367]*kernel[7]+tmp[368]*kernel[8];
				ans[268]<=tmp[167]*kernel[0]+tmp[168]*kernel[1]+tmp[169]*kernel[2]+tmp[267]*kernel[3]+tmp[268]*kernel[4]+tmp[269]*kernel[5]+tmp[367]*kernel[6]+tmp[368]*kernel[7]+tmp[369]*kernel[8];
				ans[269]<=tmp[168]*kernel[0]+tmp[169]*kernel[1]+tmp[170]*kernel[2]+tmp[268]*kernel[3]+tmp[269]*kernel[4]+tmp[270]*kernel[5]+tmp[368]*kernel[6]+tmp[369]*kernel[7]+tmp[370]*kernel[8];
				ans[270]<=tmp[169]*kernel[0]+tmp[170]*kernel[1]+tmp[171]*kernel[2]+tmp[269]*kernel[3]+tmp[270]*kernel[4]+tmp[271]*kernel[5]+tmp[369]*kernel[6]+tmp[370]*kernel[7]+tmp[371]*kernel[8];
				ans[271]<=tmp[170]*kernel[0]+tmp[171]*kernel[1]+tmp[172]*kernel[2]+tmp[270]*kernel[3]+tmp[271]*kernel[4]+tmp[272]*kernel[5]+tmp[370]*kernel[6]+tmp[371]*kernel[7]+tmp[372]*kernel[8];
				ans[272]<=tmp[171]*kernel[0]+tmp[172]*kernel[1]+tmp[173]*kernel[2]+tmp[271]*kernel[3]+tmp[272]*kernel[4]+tmp[273]*kernel[5]+tmp[371]*kernel[6]+tmp[372]*kernel[7]+tmp[373]*kernel[8];
				ans[273]<=tmp[172]*kernel[0]+tmp[173]*kernel[1]+tmp[174]*kernel[2]+tmp[272]*kernel[3]+tmp[273]*kernel[4]+tmp[274]*kernel[5]+tmp[372]*kernel[6]+tmp[373]*kernel[7]+tmp[374]*kernel[8];
				ans[274]<=tmp[173]*kernel[0]+tmp[174]*kernel[1]+tmp[175]*kernel[2]+tmp[273]*kernel[3]+tmp[274]*kernel[4]+tmp[275]*kernel[5]+tmp[373]*kernel[6]+tmp[374]*kernel[7]+tmp[375]*kernel[8];
				ans[275]<=tmp[174]*kernel[0]+tmp[175]*kernel[1]+tmp[176]*kernel[2]+tmp[274]*kernel[3]+tmp[275]*kernel[4]+tmp[276]*kernel[5]+tmp[374]*kernel[6]+tmp[375]*kernel[7]+tmp[376]*kernel[8];
				ans[276]<=tmp[175]*kernel[0]+tmp[176]*kernel[1]+tmp[177]*kernel[2]+tmp[275]*kernel[3]+tmp[276]*kernel[4]+tmp[277]*kernel[5]+tmp[375]*kernel[6]+tmp[376]*kernel[7]+tmp[377]*kernel[8];
				ans[277]<=tmp[176]*kernel[0]+tmp[177]*kernel[1]+tmp[178]*kernel[2]+tmp[276]*kernel[3]+tmp[277]*kernel[4]+tmp[278]*kernel[5]+tmp[376]*kernel[6]+tmp[377]*kernel[7]+tmp[378]*kernel[8];
				ans[278]<=tmp[177]*kernel[0]+tmp[178]*kernel[1]+tmp[179]*kernel[2]+tmp[277]*kernel[3]+tmp[278]*kernel[4]+tmp[279]*kernel[5]+tmp[377]*kernel[6]+tmp[378]*kernel[7]+tmp[379]*kernel[8];
				ans[279]<=tmp[178]*kernel[0]+tmp[179]*kernel[1]+tmp[180]*kernel[2]+tmp[278]*kernel[3]+tmp[279]*kernel[4]+tmp[280]*kernel[5]+tmp[378]*kernel[6]+tmp[379]*kernel[7]+tmp[380]*kernel[8];
				ans[280]<=tmp[179]*kernel[0]+tmp[180]*kernel[1]+tmp[181]*kernel[2]+tmp[279]*kernel[3]+tmp[280]*kernel[4]+tmp[281]*kernel[5]+tmp[379]*kernel[6]+tmp[380]*kernel[7]+tmp[381]*kernel[8];
				ans[281]<=tmp[180]*kernel[0]+tmp[181]*kernel[1]+tmp[182]*kernel[2]+tmp[280]*kernel[3]+tmp[281]*kernel[4]+tmp[282]*kernel[5]+tmp[380]*kernel[6]+tmp[381]*kernel[7]+tmp[382]*kernel[8];
				ans[282]<=tmp[181]*kernel[0]+tmp[182]*kernel[1]+tmp[183]*kernel[2]+tmp[281]*kernel[3]+tmp[282]*kernel[4]+tmp[283]*kernel[5]+tmp[381]*kernel[6]+tmp[382]*kernel[7]+tmp[383]*kernel[8];
				ans[283]<=tmp[182]*kernel[0]+tmp[183]*kernel[1]+tmp[184]*kernel[2]+tmp[282]*kernel[3]+tmp[283]*kernel[4]+tmp[284]*kernel[5]+tmp[382]*kernel[6]+tmp[383]*kernel[7]+tmp[384]*kernel[8];
				ans[284]<=tmp[183]*kernel[0]+tmp[184]*kernel[1]+tmp[185]*kernel[2]+tmp[283]*kernel[3]+tmp[284]*kernel[4]+tmp[285]*kernel[5]+tmp[383]*kernel[6]+tmp[384]*kernel[7]+tmp[385]*kernel[8];
				ans[285]<=tmp[184]*kernel[0]+tmp[185]*kernel[1]+tmp[186]*kernel[2]+tmp[284]*kernel[3]+tmp[285]*kernel[4]+tmp[286]*kernel[5]+tmp[384]*kernel[6]+tmp[385]*kernel[7]+tmp[386]*kernel[8];
				ans[286]<=tmp[185]*kernel[0]+tmp[186]*kernel[1]+tmp[187]*kernel[2]+tmp[285]*kernel[3]+tmp[286]*kernel[4]+tmp[287]*kernel[5]+tmp[385]*kernel[6]+tmp[386]*kernel[7]+tmp[387]*kernel[8];
				ans[287]<=tmp[186]*kernel[0]+tmp[187]*kernel[1]+tmp[188]*kernel[2]+tmp[286]*kernel[3]+tmp[287]*kernel[4]+tmp[288]*kernel[5]+tmp[386]*kernel[6]+tmp[387]*kernel[7]+tmp[388]*kernel[8];
				ans[288]<=tmp[187]*kernel[0]+tmp[188]*kernel[1]+tmp[189]*kernel[2]+tmp[287]*kernel[3]+tmp[288]*kernel[4]+tmp[289]*kernel[5]+tmp[387]*kernel[6]+tmp[388]*kernel[7]+tmp[389]*kernel[8];
				ans[289]<=tmp[188]*kernel[0]+tmp[189]*kernel[1]+tmp[190]*kernel[2]+tmp[288]*kernel[3]+tmp[289]*kernel[4]+tmp[290]*kernel[5]+tmp[388]*kernel[6]+tmp[389]*kernel[7]+tmp[390]*kernel[8];
				ans[290]<=tmp[189]*kernel[0]+tmp[190]*kernel[1]+tmp[191]*kernel[2]+tmp[289]*kernel[3]+tmp[290]*kernel[4]+tmp[291]*kernel[5]+tmp[389]*kernel[6]+tmp[390]*kernel[7]+tmp[391]*kernel[8];
				ans[291]<=tmp[190]*kernel[0]+tmp[191]*kernel[1]+tmp[192]*kernel[2]+tmp[290]*kernel[3]+tmp[291]*kernel[4]+tmp[292]*kernel[5]+tmp[390]*kernel[6]+tmp[391]*kernel[7]+tmp[392]*kernel[8];
				ans[292]<=tmp[191]*kernel[0]+tmp[192]*kernel[1]+tmp[193]*kernel[2]+tmp[291]*kernel[3]+tmp[292]*kernel[4]+tmp[293]*kernel[5]+tmp[391]*kernel[6]+tmp[392]*kernel[7]+tmp[393]*kernel[8];
				ans[293]<=tmp[192]*kernel[0]+tmp[193]*kernel[1]+tmp[194]*kernel[2]+tmp[292]*kernel[3]+tmp[293]*kernel[4]+tmp[294]*kernel[5]+tmp[392]*kernel[6]+tmp[393]*kernel[7]+tmp[394]*kernel[8];
				ans[294]<=tmp[193]*kernel[0]+tmp[194]*kernel[1]+tmp[195]*kernel[2]+tmp[293]*kernel[3]+tmp[294]*kernel[4]+tmp[295]*kernel[5]+tmp[393]*kernel[6]+tmp[394]*kernel[7]+tmp[395]*kernel[8];
				ans[295]<=tmp[194]*kernel[0]+tmp[195]*kernel[1]+tmp[196]*kernel[2]+tmp[294]*kernel[3]+tmp[295]*kernel[4]+tmp[296]*kernel[5]+tmp[394]*kernel[6]+tmp[395]*kernel[7]+tmp[396]*kernel[8];
				ans[296]<=tmp[195]*kernel[0]+tmp[196]*kernel[1]+tmp[197]*kernel[2]+tmp[295]*kernel[3]+tmp[296]*kernel[4]+tmp[297]*kernel[5]+tmp[395]*kernel[6]+tmp[396]*kernel[7]+tmp[397]*kernel[8];
				ans[297]<=tmp[196]*kernel[0]+tmp[197]*kernel[1]+tmp[198]*kernel[2]+tmp[296]*kernel[3]+tmp[297]*kernel[4]+tmp[298]*kernel[5]+tmp[396]*kernel[6]+tmp[397]*kernel[7]+tmp[398]*kernel[8];
				ans[298]<=tmp[197]*kernel[0]+tmp[198]*kernel[1]+tmp[199]*kernel[2]+tmp[297]*kernel[3]+tmp[298]*kernel[4]+tmp[299]*kernel[5]+tmp[397]*kernel[6]+tmp[398]*kernel[7]+tmp[399]*kernel[8];
				ans[299]<=tmp[198]*kernel[0]+tmp[199]*kernel[1]+tmp[298]*kernel[3]+tmp[299]*kernel[4]+tmp[398]*kernel[6]+tmp[399]*kernel[7];
				ans[300]<=tmp[200]*kernel[1]+tmp[201]*kernel[2]+tmp[300]*kernel[4]+tmp[301]*kernel[5]+tmp[400]*kernel[7]+tmp[401]*kernel[8];
				ans[301]<=tmp[200]*kernel[0]+tmp[201]*kernel[1]+tmp[202]*kernel[2]+tmp[300]*kernel[3]+tmp[301]*kernel[4]+tmp[302]*kernel[5]+tmp[400]*kernel[6]+tmp[401]*kernel[7]+tmp[402]*kernel[8];
				ans[302]<=tmp[201]*kernel[0]+tmp[202]*kernel[1]+tmp[203]*kernel[2]+tmp[301]*kernel[3]+tmp[302]*kernel[4]+tmp[303]*kernel[5]+tmp[401]*kernel[6]+tmp[402]*kernel[7]+tmp[403]*kernel[8];
				ans[303]<=tmp[202]*kernel[0]+tmp[203]*kernel[1]+tmp[204]*kernel[2]+tmp[302]*kernel[3]+tmp[303]*kernel[4]+tmp[304]*kernel[5]+tmp[402]*kernel[6]+tmp[403]*kernel[7]+tmp[404]*kernel[8];
				ans[304]<=tmp[203]*kernel[0]+tmp[204]*kernel[1]+tmp[205]*kernel[2]+tmp[303]*kernel[3]+tmp[304]*kernel[4]+tmp[305]*kernel[5]+tmp[403]*kernel[6]+tmp[404]*kernel[7]+tmp[405]*kernel[8];
				ans[305]<=tmp[204]*kernel[0]+tmp[205]*kernel[1]+tmp[206]*kernel[2]+tmp[304]*kernel[3]+tmp[305]*kernel[4]+tmp[306]*kernel[5]+tmp[404]*kernel[6]+tmp[405]*kernel[7]+tmp[406]*kernel[8];
				ans[306]<=tmp[205]*kernel[0]+tmp[206]*kernel[1]+tmp[207]*kernel[2]+tmp[305]*kernel[3]+tmp[306]*kernel[4]+tmp[307]*kernel[5]+tmp[405]*kernel[6]+tmp[406]*kernel[7]+tmp[407]*kernel[8];
				ans[307]<=tmp[206]*kernel[0]+tmp[207]*kernel[1]+tmp[208]*kernel[2]+tmp[306]*kernel[3]+tmp[307]*kernel[4]+tmp[308]*kernel[5]+tmp[406]*kernel[6]+tmp[407]*kernel[7]+tmp[408]*kernel[8];
				ans[308]<=tmp[207]*kernel[0]+tmp[208]*kernel[1]+tmp[209]*kernel[2]+tmp[307]*kernel[3]+tmp[308]*kernel[4]+tmp[309]*kernel[5]+tmp[407]*kernel[6]+tmp[408]*kernel[7]+tmp[409]*kernel[8];
				ans[309]<=tmp[208]*kernel[0]+tmp[209]*kernel[1]+tmp[210]*kernel[2]+tmp[308]*kernel[3]+tmp[309]*kernel[4]+tmp[310]*kernel[5]+tmp[408]*kernel[6]+tmp[409]*kernel[7]+tmp[410]*kernel[8];
				ans[310]<=tmp[209]*kernel[0]+tmp[210]*kernel[1]+tmp[211]*kernel[2]+tmp[309]*kernel[3]+tmp[310]*kernel[4]+tmp[311]*kernel[5]+tmp[409]*kernel[6]+tmp[410]*kernel[7]+tmp[411]*kernel[8];
				ans[311]<=tmp[210]*kernel[0]+tmp[211]*kernel[1]+tmp[212]*kernel[2]+tmp[310]*kernel[3]+tmp[311]*kernel[4]+tmp[312]*kernel[5]+tmp[410]*kernel[6]+tmp[411]*kernel[7]+tmp[412]*kernel[8];
				ans[312]<=tmp[211]*kernel[0]+tmp[212]*kernel[1]+tmp[213]*kernel[2]+tmp[311]*kernel[3]+tmp[312]*kernel[4]+tmp[313]*kernel[5]+tmp[411]*kernel[6]+tmp[412]*kernel[7]+tmp[413]*kernel[8];
				ans[313]<=tmp[212]*kernel[0]+tmp[213]*kernel[1]+tmp[214]*kernel[2]+tmp[312]*kernel[3]+tmp[313]*kernel[4]+tmp[314]*kernel[5]+tmp[412]*kernel[6]+tmp[413]*kernel[7]+tmp[414]*kernel[8];
				ans[314]<=tmp[213]*kernel[0]+tmp[214]*kernel[1]+tmp[215]*kernel[2]+tmp[313]*kernel[3]+tmp[314]*kernel[4]+tmp[315]*kernel[5]+tmp[413]*kernel[6]+tmp[414]*kernel[7]+tmp[415]*kernel[8];
				ans[315]<=tmp[214]*kernel[0]+tmp[215]*kernel[1]+tmp[216]*kernel[2]+tmp[314]*kernel[3]+tmp[315]*kernel[4]+tmp[316]*kernel[5]+tmp[414]*kernel[6]+tmp[415]*kernel[7]+tmp[416]*kernel[8];
				ans[316]<=tmp[215]*kernel[0]+tmp[216]*kernel[1]+tmp[217]*kernel[2]+tmp[315]*kernel[3]+tmp[316]*kernel[4]+tmp[317]*kernel[5]+tmp[415]*kernel[6]+tmp[416]*kernel[7]+tmp[417]*kernel[8];
				ans[317]<=tmp[216]*kernel[0]+tmp[217]*kernel[1]+tmp[218]*kernel[2]+tmp[316]*kernel[3]+tmp[317]*kernel[4]+tmp[318]*kernel[5]+tmp[416]*kernel[6]+tmp[417]*kernel[7]+tmp[418]*kernel[8];
				ans[318]<=tmp[217]*kernel[0]+tmp[218]*kernel[1]+tmp[219]*kernel[2]+tmp[317]*kernel[3]+tmp[318]*kernel[4]+tmp[319]*kernel[5]+tmp[417]*kernel[6]+tmp[418]*kernel[7]+tmp[419]*kernel[8];
				ans[319]<=tmp[218]*kernel[0]+tmp[219]*kernel[1]+tmp[220]*kernel[2]+tmp[318]*kernel[3]+tmp[319]*kernel[4]+tmp[320]*kernel[5]+tmp[418]*kernel[6]+tmp[419]*kernel[7]+tmp[420]*kernel[8];
				ans[320]<=tmp[219]*kernel[0]+tmp[220]*kernel[1]+tmp[221]*kernel[2]+tmp[319]*kernel[3]+tmp[320]*kernel[4]+tmp[321]*kernel[5]+tmp[419]*kernel[6]+tmp[420]*kernel[7]+tmp[421]*kernel[8];
				ans[321]<=tmp[220]*kernel[0]+tmp[221]*kernel[1]+tmp[222]*kernel[2]+tmp[320]*kernel[3]+tmp[321]*kernel[4]+tmp[322]*kernel[5]+tmp[420]*kernel[6]+tmp[421]*kernel[7]+tmp[422]*kernel[8];
				ans[322]<=tmp[221]*kernel[0]+tmp[222]*kernel[1]+tmp[223]*kernel[2]+tmp[321]*kernel[3]+tmp[322]*kernel[4]+tmp[323]*kernel[5]+tmp[421]*kernel[6]+tmp[422]*kernel[7]+tmp[423]*kernel[8];
				ans[323]<=tmp[222]*kernel[0]+tmp[223]*kernel[1]+tmp[224]*kernel[2]+tmp[322]*kernel[3]+tmp[323]*kernel[4]+tmp[324]*kernel[5]+tmp[422]*kernel[6]+tmp[423]*kernel[7]+tmp[424]*kernel[8];
				ans[324]<=tmp[223]*kernel[0]+tmp[224]*kernel[1]+tmp[225]*kernel[2]+tmp[323]*kernel[3]+tmp[324]*kernel[4]+tmp[325]*kernel[5]+tmp[423]*kernel[6]+tmp[424]*kernel[7]+tmp[425]*kernel[8];
				ans[325]<=tmp[224]*kernel[0]+tmp[225]*kernel[1]+tmp[226]*kernel[2]+tmp[324]*kernel[3]+tmp[325]*kernel[4]+tmp[326]*kernel[5]+tmp[424]*kernel[6]+tmp[425]*kernel[7]+tmp[426]*kernel[8];
				ans[326]<=tmp[225]*kernel[0]+tmp[226]*kernel[1]+tmp[227]*kernel[2]+tmp[325]*kernel[3]+tmp[326]*kernel[4]+tmp[327]*kernel[5]+tmp[425]*kernel[6]+tmp[426]*kernel[7]+tmp[427]*kernel[8];
				ans[327]<=tmp[226]*kernel[0]+tmp[227]*kernel[1]+tmp[228]*kernel[2]+tmp[326]*kernel[3]+tmp[327]*kernel[4]+tmp[328]*kernel[5]+tmp[426]*kernel[6]+tmp[427]*kernel[7]+tmp[428]*kernel[8];
				ans[328]<=tmp[227]*kernel[0]+tmp[228]*kernel[1]+tmp[229]*kernel[2]+tmp[327]*kernel[3]+tmp[328]*kernel[4]+tmp[329]*kernel[5]+tmp[427]*kernel[6]+tmp[428]*kernel[7]+tmp[429]*kernel[8];
				ans[329]<=tmp[228]*kernel[0]+tmp[229]*kernel[1]+tmp[230]*kernel[2]+tmp[328]*kernel[3]+tmp[329]*kernel[4]+tmp[330]*kernel[5]+tmp[428]*kernel[6]+tmp[429]*kernel[7]+tmp[430]*kernel[8];
				ans[330]<=tmp[229]*kernel[0]+tmp[230]*kernel[1]+tmp[231]*kernel[2]+tmp[329]*kernel[3]+tmp[330]*kernel[4]+tmp[331]*kernel[5]+tmp[429]*kernel[6]+tmp[430]*kernel[7]+tmp[431]*kernel[8];
				ans[331]<=tmp[230]*kernel[0]+tmp[231]*kernel[1]+tmp[232]*kernel[2]+tmp[330]*kernel[3]+tmp[331]*kernel[4]+tmp[332]*kernel[5]+tmp[430]*kernel[6]+tmp[431]*kernel[7]+tmp[432]*kernel[8];
				ans[332]<=tmp[231]*kernel[0]+tmp[232]*kernel[1]+tmp[233]*kernel[2]+tmp[331]*kernel[3]+tmp[332]*kernel[4]+tmp[333]*kernel[5]+tmp[431]*kernel[6]+tmp[432]*kernel[7]+tmp[433]*kernel[8];
				ans[333]<=tmp[232]*kernel[0]+tmp[233]*kernel[1]+tmp[234]*kernel[2]+tmp[332]*kernel[3]+tmp[333]*kernel[4]+tmp[334]*kernel[5]+tmp[432]*kernel[6]+tmp[433]*kernel[7]+tmp[434]*kernel[8];
				ans[334]<=tmp[233]*kernel[0]+tmp[234]*kernel[1]+tmp[235]*kernel[2]+tmp[333]*kernel[3]+tmp[334]*kernel[4]+tmp[335]*kernel[5]+tmp[433]*kernel[6]+tmp[434]*kernel[7]+tmp[435]*kernel[8];
				ans[335]<=tmp[234]*kernel[0]+tmp[235]*kernel[1]+tmp[236]*kernel[2]+tmp[334]*kernel[3]+tmp[335]*kernel[4]+tmp[336]*kernel[5]+tmp[434]*kernel[6]+tmp[435]*kernel[7]+tmp[436]*kernel[8];
				ans[336]<=tmp[235]*kernel[0]+tmp[236]*kernel[1]+tmp[237]*kernel[2]+tmp[335]*kernel[3]+tmp[336]*kernel[4]+tmp[337]*kernel[5]+tmp[435]*kernel[6]+tmp[436]*kernel[7]+tmp[437]*kernel[8];
				ans[337]<=tmp[236]*kernel[0]+tmp[237]*kernel[1]+tmp[238]*kernel[2]+tmp[336]*kernel[3]+tmp[337]*kernel[4]+tmp[338]*kernel[5]+tmp[436]*kernel[6]+tmp[437]*kernel[7]+tmp[438]*kernel[8];
				ans[338]<=tmp[237]*kernel[0]+tmp[238]*kernel[1]+tmp[239]*kernel[2]+tmp[337]*kernel[3]+tmp[338]*kernel[4]+tmp[339]*kernel[5]+tmp[437]*kernel[6]+tmp[438]*kernel[7]+tmp[439]*kernel[8];
				ans[339]<=tmp[238]*kernel[0]+tmp[239]*kernel[1]+tmp[240]*kernel[2]+tmp[338]*kernel[3]+tmp[339]*kernel[4]+tmp[340]*kernel[5]+tmp[438]*kernel[6]+tmp[439]*kernel[7]+tmp[440]*kernel[8];
				ans[340]<=tmp[239]*kernel[0]+tmp[240]*kernel[1]+tmp[241]*kernel[2]+tmp[339]*kernel[3]+tmp[340]*kernel[4]+tmp[341]*kernel[5]+tmp[439]*kernel[6]+tmp[440]*kernel[7]+tmp[441]*kernel[8];
				ans[341]<=tmp[240]*kernel[0]+tmp[241]*kernel[1]+tmp[242]*kernel[2]+tmp[340]*kernel[3]+tmp[341]*kernel[4]+tmp[342]*kernel[5]+tmp[440]*kernel[6]+tmp[441]*kernel[7]+tmp[442]*kernel[8];
				ans[342]<=tmp[241]*kernel[0]+tmp[242]*kernel[1]+tmp[243]*kernel[2]+tmp[341]*kernel[3]+tmp[342]*kernel[4]+tmp[343]*kernel[5]+tmp[441]*kernel[6]+tmp[442]*kernel[7]+tmp[443]*kernel[8];
				ans[343]<=tmp[242]*kernel[0]+tmp[243]*kernel[1]+tmp[244]*kernel[2]+tmp[342]*kernel[3]+tmp[343]*kernel[4]+tmp[344]*kernel[5]+tmp[442]*kernel[6]+tmp[443]*kernel[7]+tmp[444]*kernel[8];
				ans[344]<=tmp[243]*kernel[0]+tmp[244]*kernel[1]+tmp[245]*kernel[2]+tmp[343]*kernel[3]+tmp[344]*kernel[4]+tmp[345]*kernel[5]+tmp[443]*kernel[6]+tmp[444]*kernel[7]+tmp[445]*kernel[8];
				ans[345]<=tmp[244]*kernel[0]+tmp[245]*kernel[1]+tmp[246]*kernel[2]+tmp[344]*kernel[3]+tmp[345]*kernel[4]+tmp[346]*kernel[5]+tmp[444]*kernel[6]+tmp[445]*kernel[7]+tmp[446]*kernel[8];
				ans[346]<=tmp[245]*kernel[0]+tmp[246]*kernel[1]+tmp[247]*kernel[2]+tmp[345]*kernel[3]+tmp[346]*kernel[4]+tmp[347]*kernel[5]+tmp[445]*kernel[6]+tmp[446]*kernel[7]+tmp[447]*kernel[8];
				ans[347]<=tmp[246]*kernel[0]+tmp[247]*kernel[1]+tmp[248]*kernel[2]+tmp[346]*kernel[3]+tmp[347]*kernel[4]+tmp[348]*kernel[5]+tmp[446]*kernel[6]+tmp[447]*kernel[7]+tmp[448]*kernel[8];
				ans[348]<=tmp[247]*kernel[0]+tmp[248]*kernel[1]+tmp[249]*kernel[2]+tmp[347]*kernel[3]+tmp[348]*kernel[4]+tmp[349]*kernel[5]+tmp[447]*kernel[6]+tmp[448]*kernel[7]+tmp[449]*kernel[8];
				ans[349]<=tmp[248]*kernel[0]+tmp[249]*kernel[1]+tmp[250]*kernel[2]+tmp[348]*kernel[3]+tmp[349]*kernel[4]+tmp[350]*kernel[5]+tmp[448]*kernel[6]+tmp[449]*kernel[7]+tmp[450]*kernel[8];
				ans[350]<=tmp[249]*kernel[0]+tmp[250]*kernel[1]+tmp[251]*kernel[2]+tmp[349]*kernel[3]+tmp[350]*kernel[4]+tmp[351]*kernel[5]+tmp[449]*kernel[6]+tmp[450]*kernel[7]+tmp[451]*kernel[8];
				ans[351]<=tmp[250]*kernel[0]+tmp[251]*kernel[1]+tmp[252]*kernel[2]+tmp[350]*kernel[3]+tmp[351]*kernel[4]+tmp[352]*kernel[5]+tmp[450]*kernel[6]+tmp[451]*kernel[7]+tmp[452]*kernel[8];
				ans[352]<=tmp[251]*kernel[0]+tmp[252]*kernel[1]+tmp[253]*kernel[2]+tmp[351]*kernel[3]+tmp[352]*kernel[4]+tmp[353]*kernel[5]+tmp[451]*kernel[6]+tmp[452]*kernel[7]+tmp[453]*kernel[8];
				ans[353]<=tmp[252]*kernel[0]+tmp[253]*kernel[1]+tmp[254]*kernel[2]+tmp[352]*kernel[3]+tmp[353]*kernel[4]+tmp[354]*kernel[5]+tmp[452]*kernel[6]+tmp[453]*kernel[7]+tmp[454]*kernel[8];
				ans[354]<=tmp[253]*kernel[0]+tmp[254]*kernel[1]+tmp[255]*kernel[2]+tmp[353]*kernel[3]+tmp[354]*kernel[4]+tmp[355]*kernel[5]+tmp[453]*kernel[6]+tmp[454]*kernel[7]+tmp[455]*kernel[8];
				ans[355]<=tmp[254]*kernel[0]+tmp[255]*kernel[1]+tmp[256]*kernel[2]+tmp[354]*kernel[3]+tmp[355]*kernel[4]+tmp[356]*kernel[5]+tmp[454]*kernel[6]+tmp[455]*kernel[7]+tmp[456]*kernel[8];
				ans[356]<=tmp[255]*kernel[0]+tmp[256]*kernel[1]+tmp[257]*kernel[2]+tmp[355]*kernel[3]+tmp[356]*kernel[4]+tmp[357]*kernel[5]+tmp[455]*kernel[6]+tmp[456]*kernel[7]+tmp[457]*kernel[8];
				ans[357]<=tmp[256]*kernel[0]+tmp[257]*kernel[1]+tmp[258]*kernel[2]+tmp[356]*kernel[3]+tmp[357]*kernel[4]+tmp[358]*kernel[5]+tmp[456]*kernel[6]+tmp[457]*kernel[7]+tmp[458]*kernel[8];
				ans[358]<=tmp[257]*kernel[0]+tmp[258]*kernel[1]+tmp[259]*kernel[2]+tmp[357]*kernel[3]+tmp[358]*kernel[4]+tmp[359]*kernel[5]+tmp[457]*kernel[6]+tmp[458]*kernel[7]+tmp[459]*kernel[8];
				ans[359]<=tmp[258]*kernel[0]+tmp[259]*kernel[1]+tmp[260]*kernel[2]+tmp[358]*kernel[3]+tmp[359]*kernel[4]+tmp[360]*kernel[5]+tmp[458]*kernel[6]+tmp[459]*kernel[7]+tmp[460]*kernel[8];
				ans[360]<=tmp[259]*kernel[0]+tmp[260]*kernel[1]+tmp[261]*kernel[2]+tmp[359]*kernel[3]+tmp[360]*kernel[4]+tmp[361]*kernel[5]+tmp[459]*kernel[6]+tmp[460]*kernel[7]+tmp[461]*kernel[8];
				ans[361]<=tmp[260]*kernel[0]+tmp[261]*kernel[1]+tmp[262]*kernel[2]+tmp[360]*kernel[3]+tmp[361]*kernel[4]+tmp[362]*kernel[5]+tmp[460]*kernel[6]+tmp[461]*kernel[7]+tmp[462]*kernel[8];
				ans[362]<=tmp[261]*kernel[0]+tmp[262]*kernel[1]+tmp[263]*kernel[2]+tmp[361]*kernel[3]+tmp[362]*kernel[4]+tmp[363]*kernel[5]+tmp[461]*kernel[6]+tmp[462]*kernel[7]+tmp[463]*kernel[8];
				ans[363]<=tmp[262]*kernel[0]+tmp[263]*kernel[1]+tmp[264]*kernel[2]+tmp[362]*kernel[3]+tmp[363]*kernel[4]+tmp[364]*kernel[5]+tmp[462]*kernel[6]+tmp[463]*kernel[7]+tmp[464]*kernel[8];
				ans[364]<=tmp[263]*kernel[0]+tmp[264]*kernel[1]+tmp[265]*kernel[2]+tmp[363]*kernel[3]+tmp[364]*kernel[4]+tmp[365]*kernel[5]+tmp[463]*kernel[6]+tmp[464]*kernel[7]+tmp[465]*kernel[8];
				ans[365]<=tmp[264]*kernel[0]+tmp[265]*kernel[1]+tmp[266]*kernel[2]+tmp[364]*kernel[3]+tmp[365]*kernel[4]+tmp[366]*kernel[5]+tmp[464]*kernel[6]+tmp[465]*kernel[7]+tmp[466]*kernel[8];
				ans[366]<=tmp[265]*kernel[0]+tmp[266]*kernel[1]+tmp[267]*kernel[2]+tmp[365]*kernel[3]+tmp[366]*kernel[4]+tmp[367]*kernel[5]+tmp[465]*kernel[6]+tmp[466]*kernel[7]+tmp[467]*kernel[8];
				ans[367]<=tmp[266]*kernel[0]+tmp[267]*kernel[1]+tmp[268]*kernel[2]+tmp[366]*kernel[3]+tmp[367]*kernel[4]+tmp[368]*kernel[5]+tmp[466]*kernel[6]+tmp[467]*kernel[7]+tmp[468]*kernel[8];
				ans[368]<=tmp[267]*kernel[0]+tmp[268]*kernel[1]+tmp[269]*kernel[2]+tmp[367]*kernel[3]+tmp[368]*kernel[4]+tmp[369]*kernel[5]+tmp[467]*kernel[6]+tmp[468]*kernel[7]+tmp[469]*kernel[8];
				ans[369]<=tmp[268]*kernel[0]+tmp[269]*kernel[1]+tmp[270]*kernel[2]+tmp[368]*kernel[3]+tmp[369]*kernel[4]+tmp[370]*kernel[5]+tmp[468]*kernel[6]+tmp[469]*kernel[7]+tmp[470]*kernel[8];
				ans[370]<=tmp[269]*kernel[0]+tmp[270]*kernel[1]+tmp[271]*kernel[2]+tmp[369]*kernel[3]+tmp[370]*kernel[4]+tmp[371]*kernel[5]+tmp[469]*kernel[6]+tmp[470]*kernel[7]+tmp[471]*kernel[8];
				ans[371]<=tmp[270]*kernel[0]+tmp[271]*kernel[1]+tmp[272]*kernel[2]+tmp[370]*kernel[3]+tmp[371]*kernel[4]+tmp[372]*kernel[5]+tmp[470]*kernel[6]+tmp[471]*kernel[7]+tmp[472]*kernel[8];
				ans[372]<=tmp[271]*kernel[0]+tmp[272]*kernel[1]+tmp[273]*kernel[2]+tmp[371]*kernel[3]+tmp[372]*kernel[4]+tmp[373]*kernel[5]+tmp[471]*kernel[6]+tmp[472]*kernel[7]+tmp[473]*kernel[8];
				ans[373]<=tmp[272]*kernel[0]+tmp[273]*kernel[1]+tmp[274]*kernel[2]+tmp[372]*kernel[3]+tmp[373]*kernel[4]+tmp[374]*kernel[5]+tmp[472]*kernel[6]+tmp[473]*kernel[7]+tmp[474]*kernel[8];
				ans[374]<=tmp[273]*kernel[0]+tmp[274]*kernel[1]+tmp[275]*kernel[2]+tmp[373]*kernel[3]+tmp[374]*kernel[4]+tmp[375]*kernel[5]+tmp[473]*kernel[6]+tmp[474]*kernel[7]+tmp[475]*kernel[8];
				ans[375]<=tmp[274]*kernel[0]+tmp[275]*kernel[1]+tmp[276]*kernel[2]+tmp[374]*kernel[3]+tmp[375]*kernel[4]+tmp[376]*kernel[5]+tmp[474]*kernel[6]+tmp[475]*kernel[7]+tmp[476]*kernel[8];
				ans[376]<=tmp[275]*kernel[0]+tmp[276]*kernel[1]+tmp[277]*kernel[2]+tmp[375]*kernel[3]+tmp[376]*kernel[4]+tmp[377]*kernel[5]+tmp[475]*kernel[6]+tmp[476]*kernel[7]+tmp[477]*kernel[8];
				ans[377]<=tmp[276]*kernel[0]+tmp[277]*kernel[1]+tmp[278]*kernel[2]+tmp[376]*kernel[3]+tmp[377]*kernel[4]+tmp[378]*kernel[5]+tmp[476]*kernel[6]+tmp[477]*kernel[7]+tmp[478]*kernel[8];
				ans[378]<=tmp[277]*kernel[0]+tmp[278]*kernel[1]+tmp[279]*kernel[2]+tmp[377]*kernel[3]+tmp[378]*kernel[4]+tmp[379]*kernel[5]+tmp[477]*kernel[6]+tmp[478]*kernel[7]+tmp[479]*kernel[8];
				ans[379]<=tmp[278]*kernel[0]+tmp[279]*kernel[1]+tmp[280]*kernel[2]+tmp[378]*kernel[3]+tmp[379]*kernel[4]+tmp[380]*kernel[5]+tmp[478]*kernel[6]+tmp[479]*kernel[7]+tmp[480]*kernel[8];
				ans[380]<=tmp[279]*kernel[0]+tmp[280]*kernel[1]+tmp[281]*kernel[2]+tmp[379]*kernel[3]+tmp[380]*kernel[4]+tmp[381]*kernel[5]+tmp[479]*kernel[6]+tmp[480]*kernel[7]+tmp[481]*kernel[8];
				ans[381]<=tmp[280]*kernel[0]+tmp[281]*kernel[1]+tmp[282]*kernel[2]+tmp[380]*kernel[3]+tmp[381]*kernel[4]+tmp[382]*kernel[5]+tmp[480]*kernel[6]+tmp[481]*kernel[7]+tmp[482]*kernel[8];
				ans[382]<=tmp[281]*kernel[0]+tmp[282]*kernel[1]+tmp[283]*kernel[2]+tmp[381]*kernel[3]+tmp[382]*kernel[4]+tmp[383]*kernel[5]+tmp[481]*kernel[6]+tmp[482]*kernel[7]+tmp[483]*kernel[8];
				ans[383]<=tmp[282]*kernel[0]+tmp[283]*kernel[1]+tmp[284]*kernel[2]+tmp[382]*kernel[3]+tmp[383]*kernel[4]+tmp[384]*kernel[5]+tmp[482]*kernel[6]+tmp[483]*kernel[7]+tmp[484]*kernel[8];
				ans[384]<=tmp[283]*kernel[0]+tmp[284]*kernel[1]+tmp[285]*kernel[2]+tmp[383]*kernel[3]+tmp[384]*kernel[4]+tmp[385]*kernel[5]+tmp[483]*kernel[6]+tmp[484]*kernel[7]+tmp[485]*kernel[8];
				ans[385]<=tmp[284]*kernel[0]+tmp[285]*kernel[1]+tmp[286]*kernel[2]+tmp[384]*kernel[3]+tmp[385]*kernel[4]+tmp[386]*kernel[5]+tmp[484]*kernel[6]+tmp[485]*kernel[7]+tmp[486]*kernel[8];
				ans[386]<=tmp[285]*kernel[0]+tmp[286]*kernel[1]+tmp[287]*kernel[2]+tmp[385]*kernel[3]+tmp[386]*kernel[4]+tmp[387]*kernel[5]+tmp[485]*kernel[6]+tmp[486]*kernel[7]+tmp[487]*kernel[8];
				ans[387]<=tmp[286]*kernel[0]+tmp[287]*kernel[1]+tmp[288]*kernel[2]+tmp[386]*kernel[3]+tmp[387]*kernel[4]+tmp[388]*kernel[5]+tmp[486]*kernel[6]+tmp[487]*kernel[7]+tmp[488]*kernel[8];
				ans[388]<=tmp[287]*kernel[0]+tmp[288]*kernel[1]+tmp[289]*kernel[2]+tmp[387]*kernel[3]+tmp[388]*kernel[4]+tmp[389]*kernel[5]+tmp[487]*kernel[6]+tmp[488]*kernel[7]+tmp[489]*kernel[8];
				ans[389]<=tmp[288]*kernel[0]+tmp[289]*kernel[1]+tmp[290]*kernel[2]+tmp[388]*kernel[3]+tmp[389]*kernel[4]+tmp[390]*kernel[5]+tmp[488]*kernel[6]+tmp[489]*kernel[7]+tmp[490]*kernel[8];
				ans[390]<=tmp[289]*kernel[0]+tmp[290]*kernel[1]+tmp[291]*kernel[2]+tmp[389]*kernel[3]+tmp[390]*kernel[4]+tmp[391]*kernel[5]+tmp[489]*kernel[6]+tmp[490]*kernel[7]+tmp[491]*kernel[8];
				ans[391]<=tmp[290]*kernel[0]+tmp[291]*kernel[1]+tmp[292]*kernel[2]+tmp[390]*kernel[3]+tmp[391]*kernel[4]+tmp[392]*kernel[5]+tmp[490]*kernel[6]+tmp[491]*kernel[7]+tmp[492]*kernel[8];
				ans[392]<=tmp[291]*kernel[0]+tmp[292]*kernel[1]+tmp[293]*kernel[2]+tmp[391]*kernel[3]+tmp[392]*kernel[4]+tmp[393]*kernel[5]+tmp[491]*kernel[6]+tmp[492]*kernel[7]+tmp[493]*kernel[8];
				ans[393]<=tmp[292]*kernel[0]+tmp[293]*kernel[1]+tmp[294]*kernel[2]+tmp[392]*kernel[3]+tmp[393]*kernel[4]+tmp[394]*kernel[5]+tmp[492]*kernel[6]+tmp[493]*kernel[7]+tmp[494]*kernel[8];
				ans[394]<=tmp[293]*kernel[0]+tmp[294]*kernel[1]+tmp[295]*kernel[2]+tmp[393]*kernel[3]+tmp[394]*kernel[4]+tmp[395]*kernel[5]+tmp[493]*kernel[6]+tmp[494]*kernel[7]+tmp[495]*kernel[8];
				ans[395]<=tmp[294]*kernel[0]+tmp[295]*kernel[1]+tmp[296]*kernel[2]+tmp[394]*kernel[3]+tmp[395]*kernel[4]+tmp[396]*kernel[5]+tmp[494]*kernel[6]+tmp[495]*kernel[7]+tmp[496]*kernel[8];
				ans[396]<=tmp[295]*kernel[0]+tmp[296]*kernel[1]+tmp[297]*kernel[2]+tmp[395]*kernel[3]+tmp[396]*kernel[4]+tmp[397]*kernel[5]+tmp[495]*kernel[6]+tmp[496]*kernel[7]+tmp[497]*kernel[8];
				ans[397]<=tmp[296]*kernel[0]+tmp[297]*kernel[1]+tmp[298]*kernel[2]+tmp[396]*kernel[3]+tmp[397]*kernel[4]+tmp[398]*kernel[5]+tmp[496]*kernel[6]+tmp[497]*kernel[7]+tmp[498]*kernel[8];
				ans[398]<=tmp[297]*kernel[0]+tmp[298]*kernel[1]+tmp[299]*kernel[2]+tmp[397]*kernel[3]+tmp[398]*kernel[4]+tmp[399]*kernel[5]+tmp[497]*kernel[6]+tmp[498]*kernel[7]+tmp[499]*kernel[8];
				ans[399]<=tmp[298]*kernel[0]+tmp[299]*kernel[1]+tmp[398]*kernel[3]+tmp[399]*kernel[4]+tmp[498]*kernel[6]+tmp[499]*kernel[7];
				ans[400]<=tmp[300]*kernel[1]+tmp[301]*kernel[2]+tmp[400]*kernel[4]+tmp[401]*kernel[5]+tmp[500]*kernel[7]+tmp[501]*kernel[8];
				ans[401]<=tmp[300]*kernel[0]+tmp[301]*kernel[1]+tmp[302]*kernel[2]+tmp[400]*kernel[3]+tmp[401]*kernel[4]+tmp[402]*kernel[5]+tmp[500]*kernel[6]+tmp[501]*kernel[7]+tmp[502]*kernel[8];
				ans[402]<=tmp[301]*kernel[0]+tmp[302]*kernel[1]+tmp[303]*kernel[2]+tmp[401]*kernel[3]+tmp[402]*kernel[4]+tmp[403]*kernel[5]+tmp[501]*kernel[6]+tmp[502]*kernel[7]+tmp[503]*kernel[8];
				ans[403]<=tmp[302]*kernel[0]+tmp[303]*kernel[1]+tmp[304]*kernel[2]+tmp[402]*kernel[3]+tmp[403]*kernel[4]+tmp[404]*kernel[5]+tmp[502]*kernel[6]+tmp[503]*kernel[7]+tmp[504]*kernel[8];
				ans[404]<=tmp[303]*kernel[0]+tmp[304]*kernel[1]+tmp[305]*kernel[2]+tmp[403]*kernel[3]+tmp[404]*kernel[4]+tmp[405]*kernel[5]+tmp[503]*kernel[6]+tmp[504]*kernel[7]+tmp[505]*kernel[8];
				ans[405]<=tmp[304]*kernel[0]+tmp[305]*kernel[1]+tmp[306]*kernel[2]+tmp[404]*kernel[3]+tmp[405]*kernel[4]+tmp[406]*kernel[5]+tmp[504]*kernel[6]+tmp[505]*kernel[7]+tmp[506]*kernel[8];
				ans[406]<=tmp[305]*kernel[0]+tmp[306]*kernel[1]+tmp[307]*kernel[2]+tmp[405]*kernel[3]+tmp[406]*kernel[4]+tmp[407]*kernel[5]+tmp[505]*kernel[6]+tmp[506]*kernel[7]+tmp[507]*kernel[8];
				ans[407]<=tmp[306]*kernel[0]+tmp[307]*kernel[1]+tmp[308]*kernel[2]+tmp[406]*kernel[3]+tmp[407]*kernel[4]+tmp[408]*kernel[5]+tmp[506]*kernel[6]+tmp[507]*kernel[7]+tmp[508]*kernel[8];
				ans[408]<=tmp[307]*kernel[0]+tmp[308]*kernel[1]+tmp[309]*kernel[2]+tmp[407]*kernel[3]+tmp[408]*kernel[4]+tmp[409]*kernel[5]+tmp[507]*kernel[6]+tmp[508]*kernel[7]+tmp[509]*kernel[8];
				ans[409]<=tmp[308]*kernel[0]+tmp[309]*kernel[1]+tmp[310]*kernel[2]+tmp[408]*kernel[3]+tmp[409]*kernel[4]+tmp[410]*kernel[5]+tmp[508]*kernel[6]+tmp[509]*kernel[7]+tmp[510]*kernel[8];
				ans[410]<=tmp[309]*kernel[0]+tmp[310]*kernel[1]+tmp[311]*kernel[2]+tmp[409]*kernel[3]+tmp[410]*kernel[4]+tmp[411]*kernel[5]+tmp[509]*kernel[6]+tmp[510]*kernel[7]+tmp[511]*kernel[8];
				ans[411]<=tmp[310]*kernel[0]+tmp[311]*kernel[1]+tmp[312]*kernel[2]+tmp[410]*kernel[3]+tmp[411]*kernel[4]+tmp[412]*kernel[5]+tmp[510]*kernel[6]+tmp[511]*kernel[7]+tmp[512]*kernel[8];
				ans[412]<=tmp[311]*kernel[0]+tmp[312]*kernel[1]+tmp[313]*kernel[2]+tmp[411]*kernel[3]+tmp[412]*kernel[4]+tmp[413]*kernel[5]+tmp[511]*kernel[6]+tmp[512]*kernel[7]+tmp[513]*kernel[8];
				ans[413]<=tmp[312]*kernel[0]+tmp[313]*kernel[1]+tmp[314]*kernel[2]+tmp[412]*kernel[3]+tmp[413]*kernel[4]+tmp[414]*kernel[5]+tmp[512]*kernel[6]+tmp[513]*kernel[7]+tmp[514]*kernel[8];
				ans[414]<=tmp[313]*kernel[0]+tmp[314]*kernel[1]+tmp[315]*kernel[2]+tmp[413]*kernel[3]+tmp[414]*kernel[4]+tmp[415]*kernel[5]+tmp[513]*kernel[6]+tmp[514]*kernel[7]+tmp[515]*kernel[8];
				ans[415]<=tmp[314]*kernel[0]+tmp[315]*kernel[1]+tmp[316]*kernel[2]+tmp[414]*kernel[3]+tmp[415]*kernel[4]+tmp[416]*kernel[5]+tmp[514]*kernel[6]+tmp[515]*kernel[7]+tmp[516]*kernel[8];
				ans[416]<=tmp[315]*kernel[0]+tmp[316]*kernel[1]+tmp[317]*kernel[2]+tmp[415]*kernel[3]+tmp[416]*kernel[4]+tmp[417]*kernel[5]+tmp[515]*kernel[6]+tmp[516]*kernel[7]+tmp[517]*kernel[8];
				ans[417]<=tmp[316]*kernel[0]+tmp[317]*kernel[1]+tmp[318]*kernel[2]+tmp[416]*kernel[3]+tmp[417]*kernel[4]+tmp[418]*kernel[5]+tmp[516]*kernel[6]+tmp[517]*kernel[7]+tmp[518]*kernel[8];
				ans[418]<=tmp[317]*kernel[0]+tmp[318]*kernel[1]+tmp[319]*kernel[2]+tmp[417]*kernel[3]+tmp[418]*kernel[4]+tmp[419]*kernel[5]+tmp[517]*kernel[6]+tmp[518]*kernel[7]+tmp[519]*kernel[8];
				ans[419]<=tmp[318]*kernel[0]+tmp[319]*kernel[1]+tmp[320]*kernel[2]+tmp[418]*kernel[3]+tmp[419]*kernel[4]+tmp[420]*kernel[5]+tmp[518]*kernel[6]+tmp[519]*kernel[7]+tmp[520]*kernel[8];
				ans[420]<=tmp[319]*kernel[0]+tmp[320]*kernel[1]+tmp[321]*kernel[2]+tmp[419]*kernel[3]+tmp[420]*kernel[4]+tmp[421]*kernel[5]+tmp[519]*kernel[6]+tmp[520]*kernel[7]+tmp[521]*kernel[8];
				ans[421]<=tmp[320]*kernel[0]+tmp[321]*kernel[1]+tmp[322]*kernel[2]+tmp[420]*kernel[3]+tmp[421]*kernel[4]+tmp[422]*kernel[5]+tmp[520]*kernel[6]+tmp[521]*kernel[7]+tmp[522]*kernel[8];
				ans[422]<=tmp[321]*kernel[0]+tmp[322]*kernel[1]+tmp[323]*kernel[2]+tmp[421]*kernel[3]+tmp[422]*kernel[4]+tmp[423]*kernel[5]+tmp[521]*kernel[6]+tmp[522]*kernel[7]+tmp[523]*kernel[8];
				ans[423]<=tmp[322]*kernel[0]+tmp[323]*kernel[1]+tmp[324]*kernel[2]+tmp[422]*kernel[3]+tmp[423]*kernel[4]+tmp[424]*kernel[5]+tmp[522]*kernel[6]+tmp[523]*kernel[7]+tmp[524]*kernel[8];
				ans[424]<=tmp[323]*kernel[0]+tmp[324]*kernel[1]+tmp[325]*kernel[2]+tmp[423]*kernel[3]+tmp[424]*kernel[4]+tmp[425]*kernel[5]+tmp[523]*kernel[6]+tmp[524]*kernel[7]+tmp[525]*kernel[8];
				ans[425]<=tmp[324]*kernel[0]+tmp[325]*kernel[1]+tmp[326]*kernel[2]+tmp[424]*kernel[3]+tmp[425]*kernel[4]+tmp[426]*kernel[5]+tmp[524]*kernel[6]+tmp[525]*kernel[7]+tmp[526]*kernel[8];
				ans[426]<=tmp[325]*kernel[0]+tmp[326]*kernel[1]+tmp[327]*kernel[2]+tmp[425]*kernel[3]+tmp[426]*kernel[4]+tmp[427]*kernel[5]+tmp[525]*kernel[6]+tmp[526]*kernel[7]+tmp[527]*kernel[8];
				ans[427]<=tmp[326]*kernel[0]+tmp[327]*kernel[1]+tmp[328]*kernel[2]+tmp[426]*kernel[3]+tmp[427]*kernel[4]+tmp[428]*kernel[5]+tmp[526]*kernel[6]+tmp[527]*kernel[7]+tmp[528]*kernel[8];
				ans[428]<=tmp[327]*kernel[0]+tmp[328]*kernel[1]+tmp[329]*kernel[2]+tmp[427]*kernel[3]+tmp[428]*kernel[4]+tmp[429]*kernel[5]+tmp[527]*kernel[6]+tmp[528]*kernel[7]+tmp[529]*kernel[8];
				ans[429]<=tmp[328]*kernel[0]+tmp[329]*kernel[1]+tmp[330]*kernel[2]+tmp[428]*kernel[3]+tmp[429]*kernel[4]+tmp[430]*kernel[5]+tmp[528]*kernel[6]+tmp[529]*kernel[7]+tmp[530]*kernel[8];
				ans[430]<=tmp[329]*kernel[0]+tmp[330]*kernel[1]+tmp[331]*kernel[2]+tmp[429]*kernel[3]+tmp[430]*kernel[4]+tmp[431]*kernel[5]+tmp[529]*kernel[6]+tmp[530]*kernel[7]+tmp[531]*kernel[8];
				ans[431]<=tmp[330]*kernel[0]+tmp[331]*kernel[1]+tmp[332]*kernel[2]+tmp[430]*kernel[3]+tmp[431]*kernel[4]+tmp[432]*kernel[5]+tmp[530]*kernel[6]+tmp[531]*kernel[7]+tmp[532]*kernel[8];
				ans[432]<=tmp[331]*kernel[0]+tmp[332]*kernel[1]+tmp[333]*kernel[2]+tmp[431]*kernel[3]+tmp[432]*kernel[4]+tmp[433]*kernel[5]+tmp[531]*kernel[6]+tmp[532]*kernel[7]+tmp[533]*kernel[8];
				ans[433]<=tmp[332]*kernel[0]+tmp[333]*kernel[1]+tmp[334]*kernel[2]+tmp[432]*kernel[3]+tmp[433]*kernel[4]+tmp[434]*kernel[5]+tmp[532]*kernel[6]+tmp[533]*kernel[7]+tmp[534]*kernel[8];
				ans[434]<=tmp[333]*kernel[0]+tmp[334]*kernel[1]+tmp[335]*kernel[2]+tmp[433]*kernel[3]+tmp[434]*kernel[4]+tmp[435]*kernel[5]+tmp[533]*kernel[6]+tmp[534]*kernel[7]+tmp[535]*kernel[8];
				ans[435]<=tmp[334]*kernel[0]+tmp[335]*kernel[1]+tmp[336]*kernel[2]+tmp[434]*kernel[3]+tmp[435]*kernel[4]+tmp[436]*kernel[5]+tmp[534]*kernel[6]+tmp[535]*kernel[7]+tmp[536]*kernel[8];
				ans[436]<=tmp[335]*kernel[0]+tmp[336]*kernel[1]+tmp[337]*kernel[2]+tmp[435]*kernel[3]+tmp[436]*kernel[4]+tmp[437]*kernel[5]+tmp[535]*kernel[6]+tmp[536]*kernel[7]+tmp[537]*kernel[8];
				ans[437]<=tmp[336]*kernel[0]+tmp[337]*kernel[1]+tmp[338]*kernel[2]+tmp[436]*kernel[3]+tmp[437]*kernel[4]+tmp[438]*kernel[5]+tmp[536]*kernel[6]+tmp[537]*kernel[7]+tmp[538]*kernel[8];
				ans[438]<=tmp[337]*kernel[0]+tmp[338]*kernel[1]+tmp[339]*kernel[2]+tmp[437]*kernel[3]+tmp[438]*kernel[4]+tmp[439]*kernel[5]+tmp[537]*kernel[6]+tmp[538]*kernel[7]+tmp[539]*kernel[8];
				ans[439]<=tmp[338]*kernel[0]+tmp[339]*kernel[1]+tmp[340]*kernel[2]+tmp[438]*kernel[3]+tmp[439]*kernel[4]+tmp[440]*kernel[5]+tmp[538]*kernel[6]+tmp[539]*kernel[7]+tmp[540]*kernel[8];
				ans[440]<=tmp[339]*kernel[0]+tmp[340]*kernel[1]+tmp[341]*kernel[2]+tmp[439]*kernel[3]+tmp[440]*kernel[4]+tmp[441]*kernel[5]+tmp[539]*kernel[6]+tmp[540]*kernel[7]+tmp[541]*kernel[8];
				ans[441]<=tmp[340]*kernel[0]+tmp[341]*kernel[1]+tmp[342]*kernel[2]+tmp[440]*kernel[3]+tmp[441]*kernel[4]+tmp[442]*kernel[5]+tmp[540]*kernel[6]+tmp[541]*kernel[7]+tmp[542]*kernel[8];
				ans[442]<=tmp[341]*kernel[0]+tmp[342]*kernel[1]+tmp[343]*kernel[2]+tmp[441]*kernel[3]+tmp[442]*kernel[4]+tmp[443]*kernel[5]+tmp[541]*kernel[6]+tmp[542]*kernel[7]+tmp[543]*kernel[8];
				ans[443]<=tmp[342]*kernel[0]+tmp[343]*kernel[1]+tmp[344]*kernel[2]+tmp[442]*kernel[3]+tmp[443]*kernel[4]+tmp[444]*kernel[5]+tmp[542]*kernel[6]+tmp[543]*kernel[7]+tmp[544]*kernel[8];
				ans[444]<=tmp[343]*kernel[0]+tmp[344]*kernel[1]+tmp[345]*kernel[2]+tmp[443]*kernel[3]+tmp[444]*kernel[4]+tmp[445]*kernel[5]+tmp[543]*kernel[6]+tmp[544]*kernel[7]+tmp[545]*kernel[8];
				ans[445]<=tmp[344]*kernel[0]+tmp[345]*kernel[1]+tmp[346]*kernel[2]+tmp[444]*kernel[3]+tmp[445]*kernel[4]+tmp[446]*kernel[5]+tmp[544]*kernel[6]+tmp[545]*kernel[7]+tmp[546]*kernel[8];
				ans[446]<=tmp[345]*kernel[0]+tmp[346]*kernel[1]+tmp[347]*kernel[2]+tmp[445]*kernel[3]+tmp[446]*kernel[4]+tmp[447]*kernel[5]+tmp[545]*kernel[6]+tmp[546]*kernel[7]+tmp[547]*kernel[8];
				ans[447]<=tmp[346]*kernel[0]+tmp[347]*kernel[1]+tmp[348]*kernel[2]+tmp[446]*kernel[3]+tmp[447]*kernel[4]+tmp[448]*kernel[5]+tmp[546]*kernel[6]+tmp[547]*kernel[7]+tmp[548]*kernel[8];
				ans[448]<=tmp[347]*kernel[0]+tmp[348]*kernel[1]+tmp[349]*kernel[2]+tmp[447]*kernel[3]+tmp[448]*kernel[4]+tmp[449]*kernel[5]+tmp[547]*kernel[6]+tmp[548]*kernel[7]+tmp[549]*kernel[8];
				ans[449]<=tmp[348]*kernel[0]+tmp[349]*kernel[1]+tmp[350]*kernel[2]+tmp[448]*kernel[3]+tmp[449]*kernel[4]+tmp[450]*kernel[5]+tmp[548]*kernel[6]+tmp[549]*kernel[7]+tmp[550]*kernel[8];
				ans[450]<=tmp[349]*kernel[0]+tmp[350]*kernel[1]+tmp[351]*kernel[2]+tmp[449]*kernel[3]+tmp[450]*kernel[4]+tmp[451]*kernel[5]+tmp[549]*kernel[6]+tmp[550]*kernel[7]+tmp[551]*kernel[8];
				ans[451]<=tmp[350]*kernel[0]+tmp[351]*kernel[1]+tmp[352]*kernel[2]+tmp[450]*kernel[3]+tmp[451]*kernel[4]+tmp[452]*kernel[5]+tmp[550]*kernel[6]+tmp[551]*kernel[7]+tmp[552]*kernel[8];
				ans[452]<=tmp[351]*kernel[0]+tmp[352]*kernel[1]+tmp[353]*kernel[2]+tmp[451]*kernel[3]+tmp[452]*kernel[4]+tmp[453]*kernel[5]+tmp[551]*kernel[6]+tmp[552]*kernel[7]+tmp[553]*kernel[8];
				ans[453]<=tmp[352]*kernel[0]+tmp[353]*kernel[1]+tmp[354]*kernel[2]+tmp[452]*kernel[3]+tmp[453]*kernel[4]+tmp[454]*kernel[5]+tmp[552]*kernel[6]+tmp[553]*kernel[7]+tmp[554]*kernel[8];
				ans[454]<=tmp[353]*kernel[0]+tmp[354]*kernel[1]+tmp[355]*kernel[2]+tmp[453]*kernel[3]+tmp[454]*kernel[4]+tmp[455]*kernel[5]+tmp[553]*kernel[6]+tmp[554]*kernel[7]+tmp[555]*kernel[8];
				ans[455]<=tmp[354]*kernel[0]+tmp[355]*kernel[1]+tmp[356]*kernel[2]+tmp[454]*kernel[3]+tmp[455]*kernel[4]+tmp[456]*kernel[5]+tmp[554]*kernel[6]+tmp[555]*kernel[7]+tmp[556]*kernel[8];
				ans[456]<=tmp[355]*kernel[0]+tmp[356]*kernel[1]+tmp[357]*kernel[2]+tmp[455]*kernel[3]+tmp[456]*kernel[4]+tmp[457]*kernel[5]+tmp[555]*kernel[6]+tmp[556]*kernel[7]+tmp[557]*kernel[8];
				ans[457]<=tmp[356]*kernel[0]+tmp[357]*kernel[1]+tmp[358]*kernel[2]+tmp[456]*kernel[3]+tmp[457]*kernel[4]+tmp[458]*kernel[5]+tmp[556]*kernel[6]+tmp[557]*kernel[7]+tmp[558]*kernel[8];
				ans[458]<=tmp[357]*kernel[0]+tmp[358]*kernel[1]+tmp[359]*kernel[2]+tmp[457]*kernel[3]+tmp[458]*kernel[4]+tmp[459]*kernel[5]+tmp[557]*kernel[6]+tmp[558]*kernel[7]+tmp[559]*kernel[8];
				ans[459]<=tmp[358]*kernel[0]+tmp[359]*kernel[1]+tmp[360]*kernel[2]+tmp[458]*kernel[3]+tmp[459]*kernel[4]+tmp[460]*kernel[5]+tmp[558]*kernel[6]+tmp[559]*kernel[7]+tmp[560]*kernel[8];
				ans[460]<=tmp[359]*kernel[0]+tmp[360]*kernel[1]+tmp[361]*kernel[2]+tmp[459]*kernel[3]+tmp[460]*kernel[4]+tmp[461]*kernel[5]+tmp[559]*kernel[6]+tmp[560]*kernel[7]+tmp[561]*kernel[8];
				ans[461]<=tmp[360]*kernel[0]+tmp[361]*kernel[1]+tmp[362]*kernel[2]+tmp[460]*kernel[3]+tmp[461]*kernel[4]+tmp[462]*kernel[5]+tmp[560]*kernel[6]+tmp[561]*kernel[7]+tmp[562]*kernel[8];
				ans[462]<=tmp[361]*kernel[0]+tmp[362]*kernel[1]+tmp[363]*kernel[2]+tmp[461]*kernel[3]+tmp[462]*kernel[4]+tmp[463]*kernel[5]+tmp[561]*kernel[6]+tmp[562]*kernel[7]+tmp[563]*kernel[8];
				ans[463]<=tmp[362]*kernel[0]+tmp[363]*kernel[1]+tmp[364]*kernel[2]+tmp[462]*kernel[3]+tmp[463]*kernel[4]+tmp[464]*kernel[5]+tmp[562]*kernel[6]+tmp[563]*kernel[7]+tmp[564]*kernel[8];
				ans[464]<=tmp[363]*kernel[0]+tmp[364]*kernel[1]+tmp[365]*kernel[2]+tmp[463]*kernel[3]+tmp[464]*kernel[4]+tmp[465]*kernel[5]+tmp[563]*kernel[6]+tmp[564]*kernel[7]+tmp[565]*kernel[8];
				ans[465]<=tmp[364]*kernel[0]+tmp[365]*kernel[1]+tmp[366]*kernel[2]+tmp[464]*kernel[3]+tmp[465]*kernel[4]+tmp[466]*kernel[5]+tmp[564]*kernel[6]+tmp[565]*kernel[7]+tmp[566]*kernel[8];
				ans[466]<=tmp[365]*kernel[0]+tmp[366]*kernel[1]+tmp[367]*kernel[2]+tmp[465]*kernel[3]+tmp[466]*kernel[4]+tmp[467]*kernel[5]+tmp[565]*kernel[6]+tmp[566]*kernel[7]+tmp[567]*kernel[8];
				ans[467]<=tmp[366]*kernel[0]+tmp[367]*kernel[1]+tmp[368]*kernel[2]+tmp[466]*kernel[3]+tmp[467]*kernel[4]+tmp[468]*kernel[5]+tmp[566]*kernel[6]+tmp[567]*kernel[7]+tmp[568]*kernel[8];
				ans[468]<=tmp[367]*kernel[0]+tmp[368]*kernel[1]+tmp[369]*kernel[2]+tmp[467]*kernel[3]+tmp[468]*kernel[4]+tmp[469]*kernel[5]+tmp[567]*kernel[6]+tmp[568]*kernel[7]+tmp[569]*kernel[8];
				ans[469]<=tmp[368]*kernel[0]+tmp[369]*kernel[1]+tmp[370]*kernel[2]+tmp[468]*kernel[3]+tmp[469]*kernel[4]+tmp[470]*kernel[5]+tmp[568]*kernel[6]+tmp[569]*kernel[7]+tmp[570]*kernel[8];
				ans[470]<=tmp[369]*kernel[0]+tmp[370]*kernel[1]+tmp[371]*kernel[2]+tmp[469]*kernel[3]+tmp[470]*kernel[4]+tmp[471]*kernel[5]+tmp[569]*kernel[6]+tmp[570]*kernel[7]+tmp[571]*kernel[8];
				ans[471]<=tmp[370]*kernel[0]+tmp[371]*kernel[1]+tmp[372]*kernel[2]+tmp[470]*kernel[3]+tmp[471]*kernel[4]+tmp[472]*kernel[5]+tmp[570]*kernel[6]+tmp[571]*kernel[7]+tmp[572]*kernel[8];
				ans[472]<=tmp[371]*kernel[0]+tmp[372]*kernel[1]+tmp[373]*kernel[2]+tmp[471]*kernel[3]+tmp[472]*kernel[4]+tmp[473]*kernel[5]+tmp[571]*kernel[6]+tmp[572]*kernel[7]+tmp[573]*kernel[8];
				ans[473]<=tmp[372]*kernel[0]+tmp[373]*kernel[1]+tmp[374]*kernel[2]+tmp[472]*kernel[3]+tmp[473]*kernel[4]+tmp[474]*kernel[5]+tmp[572]*kernel[6]+tmp[573]*kernel[7]+tmp[574]*kernel[8];
				ans[474]<=tmp[373]*kernel[0]+tmp[374]*kernel[1]+tmp[375]*kernel[2]+tmp[473]*kernel[3]+tmp[474]*kernel[4]+tmp[475]*kernel[5]+tmp[573]*kernel[6]+tmp[574]*kernel[7]+tmp[575]*kernel[8];
				ans[475]<=tmp[374]*kernel[0]+tmp[375]*kernel[1]+tmp[376]*kernel[2]+tmp[474]*kernel[3]+tmp[475]*kernel[4]+tmp[476]*kernel[5]+tmp[574]*kernel[6]+tmp[575]*kernel[7]+tmp[576]*kernel[8];
				ans[476]<=tmp[375]*kernel[0]+tmp[376]*kernel[1]+tmp[377]*kernel[2]+tmp[475]*kernel[3]+tmp[476]*kernel[4]+tmp[477]*kernel[5]+tmp[575]*kernel[6]+tmp[576]*kernel[7]+tmp[577]*kernel[8];
				ans[477]<=tmp[376]*kernel[0]+tmp[377]*kernel[1]+tmp[378]*kernel[2]+tmp[476]*kernel[3]+tmp[477]*kernel[4]+tmp[478]*kernel[5]+tmp[576]*kernel[6]+tmp[577]*kernel[7]+tmp[578]*kernel[8];
				ans[478]<=tmp[377]*kernel[0]+tmp[378]*kernel[1]+tmp[379]*kernel[2]+tmp[477]*kernel[3]+tmp[478]*kernel[4]+tmp[479]*kernel[5]+tmp[577]*kernel[6]+tmp[578]*kernel[7]+tmp[579]*kernel[8];
				ans[479]<=tmp[378]*kernel[0]+tmp[379]*kernel[1]+tmp[380]*kernel[2]+tmp[478]*kernel[3]+tmp[479]*kernel[4]+tmp[480]*kernel[5]+tmp[578]*kernel[6]+tmp[579]*kernel[7]+tmp[580]*kernel[8];
				ans[480]<=tmp[379]*kernel[0]+tmp[380]*kernel[1]+tmp[381]*kernel[2]+tmp[479]*kernel[3]+tmp[480]*kernel[4]+tmp[481]*kernel[5]+tmp[579]*kernel[6]+tmp[580]*kernel[7]+tmp[581]*kernel[8];
				ans[481]<=tmp[380]*kernel[0]+tmp[381]*kernel[1]+tmp[382]*kernel[2]+tmp[480]*kernel[3]+tmp[481]*kernel[4]+tmp[482]*kernel[5]+tmp[580]*kernel[6]+tmp[581]*kernel[7]+tmp[582]*kernel[8];
				ans[482]<=tmp[381]*kernel[0]+tmp[382]*kernel[1]+tmp[383]*kernel[2]+tmp[481]*kernel[3]+tmp[482]*kernel[4]+tmp[483]*kernel[5]+tmp[581]*kernel[6]+tmp[582]*kernel[7]+tmp[583]*kernel[8];
				ans[483]<=tmp[382]*kernel[0]+tmp[383]*kernel[1]+tmp[384]*kernel[2]+tmp[482]*kernel[3]+tmp[483]*kernel[4]+tmp[484]*kernel[5]+tmp[582]*kernel[6]+tmp[583]*kernel[7]+tmp[584]*kernel[8];
				ans[484]<=tmp[383]*kernel[0]+tmp[384]*kernel[1]+tmp[385]*kernel[2]+tmp[483]*kernel[3]+tmp[484]*kernel[4]+tmp[485]*kernel[5]+tmp[583]*kernel[6]+tmp[584]*kernel[7]+tmp[585]*kernel[8];
				ans[485]<=tmp[384]*kernel[0]+tmp[385]*kernel[1]+tmp[386]*kernel[2]+tmp[484]*kernel[3]+tmp[485]*kernel[4]+tmp[486]*kernel[5]+tmp[584]*kernel[6]+tmp[585]*kernel[7]+tmp[586]*kernel[8];
				ans[486]<=tmp[385]*kernel[0]+tmp[386]*kernel[1]+tmp[387]*kernel[2]+tmp[485]*kernel[3]+tmp[486]*kernel[4]+tmp[487]*kernel[5]+tmp[585]*kernel[6]+tmp[586]*kernel[7]+tmp[587]*kernel[8];
				ans[487]<=tmp[386]*kernel[0]+tmp[387]*kernel[1]+tmp[388]*kernel[2]+tmp[486]*kernel[3]+tmp[487]*kernel[4]+tmp[488]*kernel[5]+tmp[586]*kernel[6]+tmp[587]*kernel[7]+tmp[588]*kernel[8];
				ans[488]<=tmp[387]*kernel[0]+tmp[388]*kernel[1]+tmp[389]*kernel[2]+tmp[487]*kernel[3]+tmp[488]*kernel[4]+tmp[489]*kernel[5]+tmp[587]*kernel[6]+tmp[588]*kernel[7]+tmp[589]*kernel[8];
				ans[489]<=tmp[388]*kernel[0]+tmp[389]*kernel[1]+tmp[390]*kernel[2]+tmp[488]*kernel[3]+tmp[489]*kernel[4]+tmp[490]*kernel[5]+tmp[588]*kernel[6]+tmp[589]*kernel[7]+tmp[590]*kernel[8];
				ans[490]<=tmp[389]*kernel[0]+tmp[390]*kernel[1]+tmp[391]*kernel[2]+tmp[489]*kernel[3]+tmp[490]*kernel[4]+tmp[491]*kernel[5]+tmp[589]*kernel[6]+tmp[590]*kernel[7]+tmp[591]*kernel[8];
				ans[491]<=tmp[390]*kernel[0]+tmp[391]*kernel[1]+tmp[392]*kernel[2]+tmp[490]*kernel[3]+tmp[491]*kernel[4]+tmp[492]*kernel[5]+tmp[590]*kernel[6]+tmp[591]*kernel[7]+tmp[592]*kernel[8];
				ans[492]<=tmp[391]*kernel[0]+tmp[392]*kernel[1]+tmp[393]*kernel[2]+tmp[491]*kernel[3]+tmp[492]*kernel[4]+tmp[493]*kernel[5]+tmp[591]*kernel[6]+tmp[592]*kernel[7]+tmp[593]*kernel[8];
				ans[493]<=tmp[392]*kernel[0]+tmp[393]*kernel[1]+tmp[394]*kernel[2]+tmp[492]*kernel[3]+tmp[493]*kernel[4]+tmp[494]*kernel[5]+tmp[592]*kernel[6]+tmp[593]*kernel[7]+tmp[594]*kernel[8];
				ans[494]<=tmp[393]*kernel[0]+tmp[394]*kernel[1]+tmp[395]*kernel[2]+tmp[493]*kernel[3]+tmp[494]*kernel[4]+tmp[495]*kernel[5]+tmp[593]*kernel[6]+tmp[594]*kernel[7]+tmp[595]*kernel[8];
				ans[495]<=tmp[394]*kernel[0]+tmp[395]*kernel[1]+tmp[396]*kernel[2]+tmp[494]*kernel[3]+tmp[495]*kernel[4]+tmp[496]*kernel[5]+tmp[594]*kernel[6]+tmp[595]*kernel[7]+tmp[596]*kernel[8];
				ans[496]<=tmp[395]*kernel[0]+tmp[396]*kernel[1]+tmp[397]*kernel[2]+tmp[495]*kernel[3]+tmp[496]*kernel[4]+tmp[497]*kernel[5]+tmp[595]*kernel[6]+tmp[596]*kernel[7]+tmp[597]*kernel[8];
				ans[497]<=tmp[396]*kernel[0]+tmp[397]*kernel[1]+tmp[398]*kernel[2]+tmp[496]*kernel[3]+tmp[497]*kernel[4]+tmp[498]*kernel[5]+tmp[596]*kernel[6]+tmp[597]*kernel[7]+tmp[598]*kernel[8];
				ans[498]<=tmp[397]*kernel[0]+tmp[398]*kernel[1]+tmp[399]*kernel[2]+tmp[497]*kernel[3]+tmp[498]*kernel[4]+tmp[499]*kernel[5]+tmp[597]*kernel[6]+tmp[598]*kernel[7]+tmp[599]*kernel[8];
				ans[499]<=tmp[398]*kernel[0]+tmp[399]*kernel[1]+tmp[498]*kernel[3]+tmp[499]*kernel[4]+tmp[598]*kernel[6]+tmp[599]*kernel[7];
				ans[500]<=tmp[400]*kernel[1]+tmp[401]*kernel[2]+tmp[500]*kernel[4]+tmp[501]*kernel[5]+tmp[600]*kernel[7]+tmp[601]*kernel[8];
				ans[501]<=tmp[400]*kernel[0]+tmp[401]*kernel[1]+tmp[402]*kernel[2]+tmp[500]*kernel[3]+tmp[501]*kernel[4]+tmp[502]*kernel[5]+tmp[600]*kernel[6]+tmp[601]*kernel[7]+tmp[602]*kernel[8];
				ans[502]<=tmp[401]*kernel[0]+tmp[402]*kernel[1]+tmp[403]*kernel[2]+tmp[501]*kernel[3]+tmp[502]*kernel[4]+tmp[503]*kernel[5]+tmp[601]*kernel[6]+tmp[602]*kernel[7]+tmp[603]*kernel[8];
				ans[503]<=tmp[402]*kernel[0]+tmp[403]*kernel[1]+tmp[404]*kernel[2]+tmp[502]*kernel[3]+tmp[503]*kernel[4]+tmp[504]*kernel[5]+tmp[602]*kernel[6]+tmp[603]*kernel[7]+tmp[604]*kernel[8];
				ans[504]<=tmp[403]*kernel[0]+tmp[404]*kernel[1]+tmp[405]*kernel[2]+tmp[503]*kernel[3]+tmp[504]*kernel[4]+tmp[505]*kernel[5]+tmp[603]*kernel[6]+tmp[604]*kernel[7]+tmp[605]*kernel[8];
				ans[505]<=tmp[404]*kernel[0]+tmp[405]*kernel[1]+tmp[406]*kernel[2]+tmp[504]*kernel[3]+tmp[505]*kernel[4]+tmp[506]*kernel[5]+tmp[604]*kernel[6]+tmp[605]*kernel[7]+tmp[606]*kernel[8];
				ans[506]<=tmp[405]*kernel[0]+tmp[406]*kernel[1]+tmp[407]*kernel[2]+tmp[505]*kernel[3]+tmp[506]*kernel[4]+tmp[507]*kernel[5]+tmp[605]*kernel[6]+tmp[606]*kernel[7]+tmp[607]*kernel[8];
				ans[507]<=tmp[406]*kernel[0]+tmp[407]*kernel[1]+tmp[408]*kernel[2]+tmp[506]*kernel[3]+tmp[507]*kernel[4]+tmp[508]*kernel[5]+tmp[606]*kernel[6]+tmp[607]*kernel[7]+tmp[608]*kernel[8];
				ans[508]<=tmp[407]*kernel[0]+tmp[408]*kernel[1]+tmp[409]*kernel[2]+tmp[507]*kernel[3]+tmp[508]*kernel[4]+tmp[509]*kernel[5]+tmp[607]*kernel[6]+tmp[608]*kernel[7]+tmp[609]*kernel[8];
				ans[509]<=tmp[408]*kernel[0]+tmp[409]*kernel[1]+tmp[410]*kernel[2]+tmp[508]*kernel[3]+tmp[509]*kernel[4]+tmp[510]*kernel[5]+tmp[608]*kernel[6]+tmp[609]*kernel[7]+tmp[610]*kernel[8];
				ans[510]<=tmp[409]*kernel[0]+tmp[410]*kernel[1]+tmp[411]*kernel[2]+tmp[509]*kernel[3]+tmp[510]*kernel[4]+tmp[511]*kernel[5]+tmp[609]*kernel[6]+tmp[610]*kernel[7]+tmp[611]*kernel[8];
				ans[511]<=tmp[410]*kernel[0]+tmp[411]*kernel[1]+tmp[412]*kernel[2]+tmp[510]*kernel[3]+tmp[511]*kernel[4]+tmp[512]*kernel[5]+tmp[610]*kernel[6]+tmp[611]*kernel[7]+tmp[612]*kernel[8];
				ans[512]<=tmp[411]*kernel[0]+tmp[412]*kernel[1]+tmp[413]*kernel[2]+tmp[511]*kernel[3]+tmp[512]*kernel[4]+tmp[513]*kernel[5]+tmp[611]*kernel[6]+tmp[612]*kernel[7]+tmp[613]*kernel[8];
				ans[513]<=tmp[412]*kernel[0]+tmp[413]*kernel[1]+tmp[414]*kernel[2]+tmp[512]*kernel[3]+tmp[513]*kernel[4]+tmp[514]*kernel[5]+tmp[612]*kernel[6]+tmp[613]*kernel[7]+tmp[614]*kernel[8];
				ans[514]<=tmp[413]*kernel[0]+tmp[414]*kernel[1]+tmp[415]*kernel[2]+tmp[513]*kernel[3]+tmp[514]*kernel[4]+tmp[515]*kernel[5]+tmp[613]*kernel[6]+tmp[614]*kernel[7]+tmp[615]*kernel[8];
				ans[515]<=tmp[414]*kernel[0]+tmp[415]*kernel[1]+tmp[416]*kernel[2]+tmp[514]*kernel[3]+tmp[515]*kernel[4]+tmp[516]*kernel[5]+tmp[614]*kernel[6]+tmp[615]*kernel[7]+tmp[616]*kernel[8];
				ans[516]<=tmp[415]*kernel[0]+tmp[416]*kernel[1]+tmp[417]*kernel[2]+tmp[515]*kernel[3]+tmp[516]*kernel[4]+tmp[517]*kernel[5]+tmp[615]*kernel[6]+tmp[616]*kernel[7]+tmp[617]*kernel[8];
				ans[517]<=tmp[416]*kernel[0]+tmp[417]*kernel[1]+tmp[418]*kernel[2]+tmp[516]*kernel[3]+tmp[517]*kernel[4]+tmp[518]*kernel[5]+tmp[616]*kernel[6]+tmp[617]*kernel[7]+tmp[618]*kernel[8];
				ans[518]<=tmp[417]*kernel[0]+tmp[418]*kernel[1]+tmp[419]*kernel[2]+tmp[517]*kernel[3]+tmp[518]*kernel[4]+tmp[519]*kernel[5]+tmp[617]*kernel[6]+tmp[618]*kernel[7]+tmp[619]*kernel[8];
				ans[519]<=tmp[418]*kernel[0]+tmp[419]*kernel[1]+tmp[420]*kernel[2]+tmp[518]*kernel[3]+tmp[519]*kernel[4]+tmp[520]*kernel[5]+tmp[618]*kernel[6]+tmp[619]*kernel[7]+tmp[620]*kernel[8];
				ans[520]<=tmp[419]*kernel[0]+tmp[420]*kernel[1]+tmp[421]*kernel[2]+tmp[519]*kernel[3]+tmp[520]*kernel[4]+tmp[521]*kernel[5]+tmp[619]*kernel[6]+tmp[620]*kernel[7]+tmp[621]*kernel[8];
				ans[521]<=tmp[420]*kernel[0]+tmp[421]*kernel[1]+tmp[422]*kernel[2]+tmp[520]*kernel[3]+tmp[521]*kernel[4]+tmp[522]*kernel[5]+tmp[620]*kernel[6]+tmp[621]*kernel[7]+tmp[622]*kernel[8];
				ans[522]<=tmp[421]*kernel[0]+tmp[422]*kernel[1]+tmp[423]*kernel[2]+tmp[521]*kernel[3]+tmp[522]*kernel[4]+tmp[523]*kernel[5]+tmp[621]*kernel[6]+tmp[622]*kernel[7]+tmp[623]*kernel[8];
				ans[523]<=tmp[422]*kernel[0]+tmp[423]*kernel[1]+tmp[424]*kernel[2]+tmp[522]*kernel[3]+tmp[523]*kernel[4]+tmp[524]*kernel[5]+tmp[622]*kernel[6]+tmp[623]*kernel[7]+tmp[624]*kernel[8];
				ans[524]<=tmp[423]*kernel[0]+tmp[424]*kernel[1]+tmp[425]*kernel[2]+tmp[523]*kernel[3]+tmp[524]*kernel[4]+tmp[525]*kernel[5]+tmp[623]*kernel[6]+tmp[624]*kernel[7]+tmp[625]*kernel[8];
				ans[525]<=tmp[424]*kernel[0]+tmp[425]*kernel[1]+tmp[426]*kernel[2]+tmp[524]*kernel[3]+tmp[525]*kernel[4]+tmp[526]*kernel[5]+tmp[624]*kernel[6]+tmp[625]*kernel[7]+tmp[626]*kernel[8];
				ans[526]<=tmp[425]*kernel[0]+tmp[426]*kernel[1]+tmp[427]*kernel[2]+tmp[525]*kernel[3]+tmp[526]*kernel[4]+tmp[527]*kernel[5]+tmp[625]*kernel[6]+tmp[626]*kernel[7]+tmp[627]*kernel[8];
				ans[527]<=tmp[426]*kernel[0]+tmp[427]*kernel[1]+tmp[428]*kernel[2]+tmp[526]*kernel[3]+tmp[527]*kernel[4]+tmp[528]*kernel[5]+tmp[626]*kernel[6]+tmp[627]*kernel[7]+tmp[628]*kernel[8];
				ans[528]<=tmp[427]*kernel[0]+tmp[428]*kernel[1]+tmp[429]*kernel[2]+tmp[527]*kernel[3]+tmp[528]*kernel[4]+tmp[529]*kernel[5]+tmp[627]*kernel[6]+tmp[628]*kernel[7]+tmp[629]*kernel[8];
				ans[529]<=tmp[428]*kernel[0]+tmp[429]*kernel[1]+tmp[430]*kernel[2]+tmp[528]*kernel[3]+tmp[529]*kernel[4]+tmp[530]*kernel[5]+tmp[628]*kernel[6]+tmp[629]*kernel[7]+tmp[630]*kernel[8];
				ans[530]<=tmp[429]*kernel[0]+tmp[430]*kernel[1]+tmp[431]*kernel[2]+tmp[529]*kernel[3]+tmp[530]*kernel[4]+tmp[531]*kernel[5]+tmp[629]*kernel[6]+tmp[630]*kernel[7]+tmp[631]*kernel[8];
				ans[531]<=tmp[430]*kernel[0]+tmp[431]*kernel[1]+tmp[432]*kernel[2]+tmp[530]*kernel[3]+tmp[531]*kernel[4]+tmp[532]*kernel[5]+tmp[630]*kernel[6]+tmp[631]*kernel[7]+tmp[632]*kernel[8];
				ans[532]<=tmp[431]*kernel[0]+tmp[432]*kernel[1]+tmp[433]*kernel[2]+tmp[531]*kernel[3]+tmp[532]*kernel[4]+tmp[533]*kernel[5]+tmp[631]*kernel[6]+tmp[632]*kernel[7]+tmp[633]*kernel[8];
				ans[533]<=tmp[432]*kernel[0]+tmp[433]*kernel[1]+tmp[434]*kernel[2]+tmp[532]*kernel[3]+tmp[533]*kernel[4]+tmp[534]*kernel[5]+tmp[632]*kernel[6]+tmp[633]*kernel[7]+tmp[634]*kernel[8];
				ans[534]<=tmp[433]*kernel[0]+tmp[434]*kernel[1]+tmp[435]*kernel[2]+tmp[533]*kernel[3]+tmp[534]*kernel[4]+tmp[535]*kernel[5]+tmp[633]*kernel[6]+tmp[634]*kernel[7]+tmp[635]*kernel[8];
				ans[535]<=tmp[434]*kernel[0]+tmp[435]*kernel[1]+tmp[436]*kernel[2]+tmp[534]*kernel[3]+tmp[535]*kernel[4]+tmp[536]*kernel[5]+tmp[634]*kernel[6]+tmp[635]*kernel[7]+tmp[636]*kernel[8];
				ans[536]<=tmp[435]*kernel[0]+tmp[436]*kernel[1]+tmp[437]*kernel[2]+tmp[535]*kernel[3]+tmp[536]*kernel[4]+tmp[537]*kernel[5]+tmp[635]*kernel[6]+tmp[636]*kernel[7]+tmp[637]*kernel[8];
				ans[537]<=tmp[436]*kernel[0]+tmp[437]*kernel[1]+tmp[438]*kernel[2]+tmp[536]*kernel[3]+tmp[537]*kernel[4]+tmp[538]*kernel[5]+tmp[636]*kernel[6]+tmp[637]*kernel[7]+tmp[638]*kernel[8];
				ans[538]<=tmp[437]*kernel[0]+tmp[438]*kernel[1]+tmp[439]*kernel[2]+tmp[537]*kernel[3]+tmp[538]*kernel[4]+tmp[539]*kernel[5]+tmp[637]*kernel[6]+tmp[638]*kernel[7]+tmp[639]*kernel[8];
				ans[539]<=tmp[438]*kernel[0]+tmp[439]*kernel[1]+tmp[440]*kernel[2]+tmp[538]*kernel[3]+tmp[539]*kernel[4]+tmp[540]*kernel[5]+tmp[638]*kernel[6]+tmp[639]*kernel[7]+tmp[640]*kernel[8];
				ans[540]<=tmp[439]*kernel[0]+tmp[440]*kernel[1]+tmp[441]*kernel[2]+tmp[539]*kernel[3]+tmp[540]*kernel[4]+tmp[541]*kernel[5]+tmp[639]*kernel[6]+tmp[640]*kernel[7]+tmp[641]*kernel[8];
				ans[541]<=tmp[440]*kernel[0]+tmp[441]*kernel[1]+tmp[442]*kernel[2]+tmp[540]*kernel[3]+tmp[541]*kernel[4]+tmp[542]*kernel[5]+tmp[640]*kernel[6]+tmp[641]*kernel[7]+tmp[642]*kernel[8];
				ans[542]<=tmp[441]*kernel[0]+tmp[442]*kernel[1]+tmp[443]*kernel[2]+tmp[541]*kernel[3]+tmp[542]*kernel[4]+tmp[543]*kernel[5]+tmp[641]*kernel[6]+tmp[642]*kernel[7]+tmp[643]*kernel[8];
				ans[543]<=tmp[442]*kernel[0]+tmp[443]*kernel[1]+tmp[444]*kernel[2]+tmp[542]*kernel[3]+tmp[543]*kernel[4]+tmp[544]*kernel[5]+tmp[642]*kernel[6]+tmp[643]*kernel[7]+tmp[644]*kernel[8];
				ans[544]<=tmp[443]*kernel[0]+tmp[444]*kernel[1]+tmp[445]*kernel[2]+tmp[543]*kernel[3]+tmp[544]*kernel[4]+tmp[545]*kernel[5]+tmp[643]*kernel[6]+tmp[644]*kernel[7]+tmp[645]*kernel[8];
				ans[545]<=tmp[444]*kernel[0]+tmp[445]*kernel[1]+tmp[446]*kernel[2]+tmp[544]*kernel[3]+tmp[545]*kernel[4]+tmp[546]*kernel[5]+tmp[644]*kernel[6]+tmp[645]*kernel[7]+tmp[646]*kernel[8];
				ans[546]<=tmp[445]*kernel[0]+tmp[446]*kernel[1]+tmp[447]*kernel[2]+tmp[545]*kernel[3]+tmp[546]*kernel[4]+tmp[547]*kernel[5]+tmp[645]*kernel[6]+tmp[646]*kernel[7]+tmp[647]*kernel[8];
				ans[547]<=tmp[446]*kernel[0]+tmp[447]*kernel[1]+tmp[448]*kernel[2]+tmp[546]*kernel[3]+tmp[547]*kernel[4]+tmp[548]*kernel[5]+tmp[646]*kernel[6]+tmp[647]*kernel[7]+tmp[648]*kernel[8];
				ans[548]<=tmp[447]*kernel[0]+tmp[448]*kernel[1]+tmp[449]*kernel[2]+tmp[547]*kernel[3]+tmp[548]*kernel[4]+tmp[549]*kernel[5]+tmp[647]*kernel[6]+tmp[648]*kernel[7]+tmp[649]*kernel[8];
				ans[549]<=tmp[448]*kernel[0]+tmp[449]*kernel[1]+tmp[450]*kernel[2]+tmp[548]*kernel[3]+tmp[549]*kernel[4]+tmp[550]*kernel[5]+tmp[648]*kernel[6]+tmp[649]*kernel[7]+tmp[650]*kernel[8];
				ans[550]<=tmp[449]*kernel[0]+tmp[450]*kernel[1]+tmp[451]*kernel[2]+tmp[549]*kernel[3]+tmp[550]*kernel[4]+tmp[551]*kernel[5]+tmp[649]*kernel[6]+tmp[650]*kernel[7]+tmp[651]*kernel[8];
				ans[551]<=tmp[450]*kernel[0]+tmp[451]*kernel[1]+tmp[452]*kernel[2]+tmp[550]*kernel[3]+tmp[551]*kernel[4]+tmp[552]*kernel[5]+tmp[650]*kernel[6]+tmp[651]*kernel[7]+tmp[652]*kernel[8];
				ans[552]<=tmp[451]*kernel[0]+tmp[452]*kernel[1]+tmp[453]*kernel[2]+tmp[551]*kernel[3]+tmp[552]*kernel[4]+tmp[553]*kernel[5]+tmp[651]*kernel[6]+tmp[652]*kernel[7]+tmp[653]*kernel[8];
				ans[553]<=tmp[452]*kernel[0]+tmp[453]*kernel[1]+tmp[454]*kernel[2]+tmp[552]*kernel[3]+tmp[553]*kernel[4]+tmp[554]*kernel[5]+tmp[652]*kernel[6]+tmp[653]*kernel[7]+tmp[654]*kernel[8];
				ans[554]<=tmp[453]*kernel[0]+tmp[454]*kernel[1]+tmp[455]*kernel[2]+tmp[553]*kernel[3]+tmp[554]*kernel[4]+tmp[555]*kernel[5]+tmp[653]*kernel[6]+tmp[654]*kernel[7]+tmp[655]*kernel[8];
				ans[555]<=tmp[454]*kernel[0]+tmp[455]*kernel[1]+tmp[456]*kernel[2]+tmp[554]*kernel[3]+tmp[555]*kernel[4]+tmp[556]*kernel[5]+tmp[654]*kernel[6]+tmp[655]*kernel[7]+tmp[656]*kernel[8];
				ans[556]<=tmp[455]*kernel[0]+tmp[456]*kernel[1]+tmp[457]*kernel[2]+tmp[555]*kernel[3]+tmp[556]*kernel[4]+tmp[557]*kernel[5]+tmp[655]*kernel[6]+tmp[656]*kernel[7]+tmp[657]*kernel[8];
				ans[557]<=tmp[456]*kernel[0]+tmp[457]*kernel[1]+tmp[458]*kernel[2]+tmp[556]*kernel[3]+tmp[557]*kernel[4]+tmp[558]*kernel[5]+tmp[656]*kernel[6]+tmp[657]*kernel[7]+tmp[658]*kernel[8];
				ans[558]<=tmp[457]*kernel[0]+tmp[458]*kernel[1]+tmp[459]*kernel[2]+tmp[557]*kernel[3]+tmp[558]*kernel[4]+tmp[559]*kernel[5]+tmp[657]*kernel[6]+tmp[658]*kernel[7]+tmp[659]*kernel[8];
				ans[559]<=tmp[458]*kernel[0]+tmp[459]*kernel[1]+tmp[460]*kernel[2]+tmp[558]*kernel[3]+tmp[559]*kernel[4]+tmp[560]*kernel[5]+tmp[658]*kernel[6]+tmp[659]*kernel[7]+tmp[660]*kernel[8];
				ans[560]<=tmp[459]*kernel[0]+tmp[460]*kernel[1]+tmp[461]*kernel[2]+tmp[559]*kernel[3]+tmp[560]*kernel[4]+tmp[561]*kernel[5]+tmp[659]*kernel[6]+tmp[660]*kernel[7]+tmp[661]*kernel[8];
				ans[561]<=tmp[460]*kernel[0]+tmp[461]*kernel[1]+tmp[462]*kernel[2]+tmp[560]*kernel[3]+tmp[561]*kernel[4]+tmp[562]*kernel[5]+tmp[660]*kernel[6]+tmp[661]*kernel[7]+tmp[662]*kernel[8];
				ans[562]<=tmp[461]*kernel[0]+tmp[462]*kernel[1]+tmp[463]*kernel[2]+tmp[561]*kernel[3]+tmp[562]*kernel[4]+tmp[563]*kernel[5]+tmp[661]*kernel[6]+tmp[662]*kernel[7]+tmp[663]*kernel[8];
				ans[563]<=tmp[462]*kernel[0]+tmp[463]*kernel[1]+tmp[464]*kernel[2]+tmp[562]*kernel[3]+tmp[563]*kernel[4]+tmp[564]*kernel[5]+tmp[662]*kernel[6]+tmp[663]*kernel[7]+tmp[664]*kernel[8];
				ans[564]<=tmp[463]*kernel[0]+tmp[464]*kernel[1]+tmp[465]*kernel[2]+tmp[563]*kernel[3]+tmp[564]*kernel[4]+tmp[565]*kernel[5]+tmp[663]*kernel[6]+tmp[664]*kernel[7]+tmp[665]*kernel[8];
				ans[565]<=tmp[464]*kernel[0]+tmp[465]*kernel[1]+tmp[466]*kernel[2]+tmp[564]*kernel[3]+tmp[565]*kernel[4]+tmp[566]*kernel[5]+tmp[664]*kernel[6]+tmp[665]*kernel[7]+tmp[666]*kernel[8];
				ans[566]<=tmp[465]*kernel[0]+tmp[466]*kernel[1]+tmp[467]*kernel[2]+tmp[565]*kernel[3]+tmp[566]*kernel[4]+tmp[567]*kernel[5]+tmp[665]*kernel[6]+tmp[666]*kernel[7]+tmp[667]*kernel[8];
				ans[567]<=tmp[466]*kernel[0]+tmp[467]*kernel[1]+tmp[468]*kernel[2]+tmp[566]*kernel[3]+tmp[567]*kernel[4]+tmp[568]*kernel[5]+tmp[666]*kernel[6]+tmp[667]*kernel[7]+tmp[668]*kernel[8];
				ans[568]<=tmp[467]*kernel[0]+tmp[468]*kernel[1]+tmp[469]*kernel[2]+tmp[567]*kernel[3]+tmp[568]*kernel[4]+tmp[569]*kernel[5]+tmp[667]*kernel[6]+tmp[668]*kernel[7]+tmp[669]*kernel[8];
				ans[569]<=tmp[468]*kernel[0]+tmp[469]*kernel[1]+tmp[470]*kernel[2]+tmp[568]*kernel[3]+tmp[569]*kernel[4]+tmp[570]*kernel[5]+tmp[668]*kernel[6]+tmp[669]*kernel[7]+tmp[670]*kernel[8];
				ans[570]<=tmp[469]*kernel[0]+tmp[470]*kernel[1]+tmp[471]*kernel[2]+tmp[569]*kernel[3]+tmp[570]*kernel[4]+tmp[571]*kernel[5]+tmp[669]*kernel[6]+tmp[670]*kernel[7]+tmp[671]*kernel[8];
				ans[571]<=tmp[470]*kernel[0]+tmp[471]*kernel[1]+tmp[472]*kernel[2]+tmp[570]*kernel[3]+tmp[571]*kernel[4]+tmp[572]*kernel[5]+tmp[670]*kernel[6]+tmp[671]*kernel[7]+tmp[672]*kernel[8];
				ans[572]<=tmp[471]*kernel[0]+tmp[472]*kernel[1]+tmp[473]*kernel[2]+tmp[571]*kernel[3]+tmp[572]*kernel[4]+tmp[573]*kernel[5]+tmp[671]*kernel[6]+tmp[672]*kernel[7]+tmp[673]*kernel[8];
				ans[573]<=tmp[472]*kernel[0]+tmp[473]*kernel[1]+tmp[474]*kernel[2]+tmp[572]*kernel[3]+tmp[573]*kernel[4]+tmp[574]*kernel[5]+tmp[672]*kernel[6]+tmp[673]*kernel[7]+tmp[674]*kernel[8];
				ans[574]<=tmp[473]*kernel[0]+tmp[474]*kernel[1]+tmp[475]*kernel[2]+tmp[573]*kernel[3]+tmp[574]*kernel[4]+tmp[575]*kernel[5]+tmp[673]*kernel[6]+tmp[674]*kernel[7]+tmp[675]*kernel[8];
				ans[575]<=tmp[474]*kernel[0]+tmp[475]*kernel[1]+tmp[476]*kernel[2]+tmp[574]*kernel[3]+tmp[575]*kernel[4]+tmp[576]*kernel[5]+tmp[674]*kernel[6]+tmp[675]*kernel[7]+tmp[676]*kernel[8];
				ans[576]<=tmp[475]*kernel[0]+tmp[476]*kernel[1]+tmp[477]*kernel[2]+tmp[575]*kernel[3]+tmp[576]*kernel[4]+tmp[577]*kernel[5]+tmp[675]*kernel[6]+tmp[676]*kernel[7]+tmp[677]*kernel[8];
				ans[577]<=tmp[476]*kernel[0]+tmp[477]*kernel[1]+tmp[478]*kernel[2]+tmp[576]*kernel[3]+tmp[577]*kernel[4]+tmp[578]*kernel[5]+tmp[676]*kernel[6]+tmp[677]*kernel[7]+tmp[678]*kernel[8];
				ans[578]<=tmp[477]*kernel[0]+tmp[478]*kernel[1]+tmp[479]*kernel[2]+tmp[577]*kernel[3]+tmp[578]*kernel[4]+tmp[579]*kernel[5]+tmp[677]*kernel[6]+tmp[678]*kernel[7]+tmp[679]*kernel[8];
				ans[579]<=tmp[478]*kernel[0]+tmp[479]*kernel[1]+tmp[480]*kernel[2]+tmp[578]*kernel[3]+tmp[579]*kernel[4]+tmp[580]*kernel[5]+tmp[678]*kernel[6]+tmp[679]*kernel[7]+tmp[680]*kernel[8];
				ans[580]<=tmp[479]*kernel[0]+tmp[480]*kernel[1]+tmp[481]*kernel[2]+tmp[579]*kernel[3]+tmp[580]*kernel[4]+tmp[581]*kernel[5]+tmp[679]*kernel[6]+tmp[680]*kernel[7]+tmp[681]*kernel[8];
				ans[581]<=tmp[480]*kernel[0]+tmp[481]*kernel[1]+tmp[482]*kernel[2]+tmp[580]*kernel[3]+tmp[581]*kernel[4]+tmp[582]*kernel[5]+tmp[680]*kernel[6]+tmp[681]*kernel[7]+tmp[682]*kernel[8];
				ans[582]<=tmp[481]*kernel[0]+tmp[482]*kernel[1]+tmp[483]*kernel[2]+tmp[581]*kernel[3]+tmp[582]*kernel[4]+tmp[583]*kernel[5]+tmp[681]*kernel[6]+tmp[682]*kernel[7]+tmp[683]*kernel[8];
				ans[583]<=tmp[482]*kernel[0]+tmp[483]*kernel[1]+tmp[484]*kernel[2]+tmp[582]*kernel[3]+tmp[583]*kernel[4]+tmp[584]*kernel[5]+tmp[682]*kernel[6]+tmp[683]*kernel[7]+tmp[684]*kernel[8];
				ans[584]<=tmp[483]*kernel[0]+tmp[484]*kernel[1]+tmp[485]*kernel[2]+tmp[583]*kernel[3]+tmp[584]*kernel[4]+tmp[585]*kernel[5]+tmp[683]*kernel[6]+tmp[684]*kernel[7]+tmp[685]*kernel[8];
				ans[585]<=tmp[484]*kernel[0]+tmp[485]*kernel[1]+tmp[486]*kernel[2]+tmp[584]*kernel[3]+tmp[585]*kernel[4]+tmp[586]*kernel[5]+tmp[684]*kernel[6]+tmp[685]*kernel[7]+tmp[686]*kernel[8];
				ans[586]<=tmp[485]*kernel[0]+tmp[486]*kernel[1]+tmp[487]*kernel[2]+tmp[585]*kernel[3]+tmp[586]*kernel[4]+tmp[587]*kernel[5]+tmp[685]*kernel[6]+tmp[686]*kernel[7]+tmp[687]*kernel[8];
				ans[587]<=tmp[486]*kernel[0]+tmp[487]*kernel[1]+tmp[488]*kernel[2]+tmp[586]*kernel[3]+tmp[587]*kernel[4]+tmp[588]*kernel[5]+tmp[686]*kernel[6]+tmp[687]*kernel[7]+tmp[688]*kernel[8];
				ans[588]<=tmp[487]*kernel[0]+tmp[488]*kernel[1]+tmp[489]*kernel[2]+tmp[587]*kernel[3]+tmp[588]*kernel[4]+tmp[589]*kernel[5]+tmp[687]*kernel[6]+tmp[688]*kernel[7]+tmp[689]*kernel[8];
				ans[589]<=tmp[488]*kernel[0]+tmp[489]*kernel[1]+tmp[490]*kernel[2]+tmp[588]*kernel[3]+tmp[589]*kernel[4]+tmp[590]*kernel[5]+tmp[688]*kernel[6]+tmp[689]*kernel[7]+tmp[690]*kernel[8];
				ans[590]<=tmp[489]*kernel[0]+tmp[490]*kernel[1]+tmp[491]*kernel[2]+tmp[589]*kernel[3]+tmp[590]*kernel[4]+tmp[591]*kernel[5]+tmp[689]*kernel[6]+tmp[690]*kernel[7]+tmp[691]*kernel[8];
				ans[591]<=tmp[490]*kernel[0]+tmp[491]*kernel[1]+tmp[492]*kernel[2]+tmp[590]*kernel[3]+tmp[591]*kernel[4]+tmp[592]*kernel[5]+tmp[690]*kernel[6]+tmp[691]*kernel[7]+tmp[692]*kernel[8];
				ans[592]<=tmp[491]*kernel[0]+tmp[492]*kernel[1]+tmp[493]*kernel[2]+tmp[591]*kernel[3]+tmp[592]*kernel[4]+tmp[593]*kernel[5]+tmp[691]*kernel[6]+tmp[692]*kernel[7]+tmp[693]*kernel[8];
				ans[593]<=tmp[492]*kernel[0]+tmp[493]*kernel[1]+tmp[494]*kernel[2]+tmp[592]*kernel[3]+tmp[593]*kernel[4]+tmp[594]*kernel[5]+tmp[692]*kernel[6]+tmp[693]*kernel[7]+tmp[694]*kernel[8];
				ans[594]<=tmp[493]*kernel[0]+tmp[494]*kernel[1]+tmp[495]*kernel[2]+tmp[593]*kernel[3]+tmp[594]*kernel[4]+tmp[595]*kernel[5]+tmp[693]*kernel[6]+tmp[694]*kernel[7]+tmp[695]*kernel[8];
				ans[595]<=tmp[494]*kernel[0]+tmp[495]*kernel[1]+tmp[496]*kernel[2]+tmp[594]*kernel[3]+tmp[595]*kernel[4]+tmp[596]*kernel[5]+tmp[694]*kernel[6]+tmp[695]*kernel[7]+tmp[696]*kernel[8];
				ans[596]<=tmp[495]*kernel[0]+tmp[496]*kernel[1]+tmp[497]*kernel[2]+tmp[595]*kernel[3]+tmp[596]*kernel[4]+tmp[597]*kernel[5]+tmp[695]*kernel[6]+tmp[696]*kernel[7]+tmp[697]*kernel[8];
				ans[597]<=tmp[496]*kernel[0]+tmp[497]*kernel[1]+tmp[498]*kernel[2]+tmp[596]*kernel[3]+tmp[597]*kernel[4]+tmp[598]*kernel[5]+tmp[696]*kernel[6]+tmp[697]*kernel[7]+tmp[698]*kernel[8];
				ans[598]<=tmp[497]*kernel[0]+tmp[498]*kernel[1]+tmp[499]*kernel[2]+tmp[597]*kernel[3]+tmp[598]*kernel[4]+tmp[599]*kernel[5]+tmp[697]*kernel[6]+tmp[698]*kernel[7]+tmp[699]*kernel[8];
				ans[599]<=tmp[498]*kernel[0]+tmp[499]*kernel[1]+tmp[598]*kernel[3]+tmp[599]*kernel[4]+tmp[698]*kernel[6]+tmp[699]*kernel[7];
				ans[600]<=tmp[500]*kernel[1]+tmp[501]*kernel[2]+tmp[600]*kernel[4]+tmp[601]*kernel[5]+tmp[700]*kernel[7]+tmp[701]*kernel[8];
				ans[601]<=tmp[500]*kernel[0]+tmp[501]*kernel[1]+tmp[502]*kernel[2]+tmp[600]*kernel[3]+tmp[601]*kernel[4]+tmp[602]*kernel[5]+tmp[700]*kernel[6]+tmp[701]*kernel[7]+tmp[702]*kernel[8];
				ans[602]<=tmp[501]*kernel[0]+tmp[502]*kernel[1]+tmp[503]*kernel[2]+tmp[601]*kernel[3]+tmp[602]*kernel[4]+tmp[603]*kernel[5]+tmp[701]*kernel[6]+tmp[702]*kernel[7]+tmp[703]*kernel[8];
				ans[603]<=tmp[502]*kernel[0]+tmp[503]*kernel[1]+tmp[504]*kernel[2]+tmp[602]*kernel[3]+tmp[603]*kernel[4]+tmp[604]*kernel[5]+tmp[702]*kernel[6]+tmp[703]*kernel[7]+tmp[704]*kernel[8];
				ans[604]<=tmp[503]*kernel[0]+tmp[504]*kernel[1]+tmp[505]*kernel[2]+tmp[603]*kernel[3]+tmp[604]*kernel[4]+tmp[605]*kernel[5]+tmp[703]*kernel[6]+tmp[704]*kernel[7]+tmp[705]*kernel[8];
				ans[605]<=tmp[504]*kernel[0]+tmp[505]*kernel[1]+tmp[506]*kernel[2]+tmp[604]*kernel[3]+tmp[605]*kernel[4]+tmp[606]*kernel[5]+tmp[704]*kernel[6]+tmp[705]*kernel[7]+tmp[706]*kernel[8];
				ans[606]<=tmp[505]*kernel[0]+tmp[506]*kernel[1]+tmp[507]*kernel[2]+tmp[605]*kernel[3]+tmp[606]*kernel[4]+tmp[607]*kernel[5]+tmp[705]*kernel[6]+tmp[706]*kernel[7]+tmp[707]*kernel[8];
				ans[607]<=tmp[506]*kernel[0]+tmp[507]*kernel[1]+tmp[508]*kernel[2]+tmp[606]*kernel[3]+tmp[607]*kernel[4]+tmp[608]*kernel[5]+tmp[706]*kernel[6]+tmp[707]*kernel[7]+tmp[708]*kernel[8];
				ans[608]<=tmp[507]*kernel[0]+tmp[508]*kernel[1]+tmp[509]*kernel[2]+tmp[607]*kernel[3]+tmp[608]*kernel[4]+tmp[609]*kernel[5]+tmp[707]*kernel[6]+tmp[708]*kernel[7]+tmp[709]*kernel[8];
				ans[609]<=tmp[508]*kernel[0]+tmp[509]*kernel[1]+tmp[510]*kernel[2]+tmp[608]*kernel[3]+tmp[609]*kernel[4]+tmp[610]*kernel[5]+tmp[708]*kernel[6]+tmp[709]*kernel[7]+tmp[710]*kernel[8];
				ans[610]<=tmp[509]*kernel[0]+tmp[510]*kernel[1]+tmp[511]*kernel[2]+tmp[609]*kernel[3]+tmp[610]*kernel[4]+tmp[611]*kernel[5]+tmp[709]*kernel[6]+tmp[710]*kernel[7]+tmp[711]*kernel[8];
				ans[611]<=tmp[510]*kernel[0]+tmp[511]*kernel[1]+tmp[512]*kernel[2]+tmp[610]*kernel[3]+tmp[611]*kernel[4]+tmp[612]*kernel[5]+tmp[710]*kernel[6]+tmp[711]*kernel[7]+tmp[712]*kernel[8];
				ans[612]<=tmp[511]*kernel[0]+tmp[512]*kernel[1]+tmp[513]*kernel[2]+tmp[611]*kernel[3]+tmp[612]*kernel[4]+tmp[613]*kernel[5]+tmp[711]*kernel[6]+tmp[712]*kernel[7]+tmp[713]*kernel[8];
				ans[613]<=tmp[512]*kernel[0]+tmp[513]*kernel[1]+tmp[514]*kernel[2]+tmp[612]*kernel[3]+tmp[613]*kernel[4]+tmp[614]*kernel[5]+tmp[712]*kernel[6]+tmp[713]*kernel[7]+tmp[714]*kernel[8];
				ans[614]<=tmp[513]*kernel[0]+tmp[514]*kernel[1]+tmp[515]*kernel[2]+tmp[613]*kernel[3]+tmp[614]*kernel[4]+tmp[615]*kernel[5]+tmp[713]*kernel[6]+tmp[714]*kernel[7]+tmp[715]*kernel[8];
				ans[615]<=tmp[514]*kernel[0]+tmp[515]*kernel[1]+tmp[516]*kernel[2]+tmp[614]*kernel[3]+tmp[615]*kernel[4]+tmp[616]*kernel[5]+tmp[714]*kernel[6]+tmp[715]*kernel[7]+tmp[716]*kernel[8];
				ans[616]<=tmp[515]*kernel[0]+tmp[516]*kernel[1]+tmp[517]*kernel[2]+tmp[615]*kernel[3]+tmp[616]*kernel[4]+tmp[617]*kernel[5]+tmp[715]*kernel[6]+tmp[716]*kernel[7]+tmp[717]*kernel[8];
				ans[617]<=tmp[516]*kernel[0]+tmp[517]*kernel[1]+tmp[518]*kernel[2]+tmp[616]*kernel[3]+tmp[617]*kernel[4]+tmp[618]*kernel[5]+tmp[716]*kernel[6]+tmp[717]*kernel[7]+tmp[718]*kernel[8];
				ans[618]<=tmp[517]*kernel[0]+tmp[518]*kernel[1]+tmp[519]*kernel[2]+tmp[617]*kernel[3]+tmp[618]*kernel[4]+tmp[619]*kernel[5]+tmp[717]*kernel[6]+tmp[718]*kernel[7]+tmp[719]*kernel[8];
				ans[619]<=tmp[518]*kernel[0]+tmp[519]*kernel[1]+tmp[520]*kernel[2]+tmp[618]*kernel[3]+tmp[619]*kernel[4]+tmp[620]*kernel[5]+tmp[718]*kernel[6]+tmp[719]*kernel[7]+tmp[720]*kernel[8];
				ans[620]<=tmp[519]*kernel[0]+tmp[520]*kernel[1]+tmp[521]*kernel[2]+tmp[619]*kernel[3]+tmp[620]*kernel[4]+tmp[621]*kernel[5]+tmp[719]*kernel[6]+tmp[720]*kernel[7]+tmp[721]*kernel[8];
				ans[621]<=tmp[520]*kernel[0]+tmp[521]*kernel[1]+tmp[522]*kernel[2]+tmp[620]*kernel[3]+tmp[621]*kernel[4]+tmp[622]*kernel[5]+tmp[720]*kernel[6]+tmp[721]*kernel[7]+tmp[722]*kernel[8];
				ans[622]<=tmp[521]*kernel[0]+tmp[522]*kernel[1]+tmp[523]*kernel[2]+tmp[621]*kernel[3]+tmp[622]*kernel[4]+tmp[623]*kernel[5]+tmp[721]*kernel[6]+tmp[722]*kernel[7]+tmp[723]*kernel[8];
				ans[623]<=tmp[522]*kernel[0]+tmp[523]*kernel[1]+tmp[524]*kernel[2]+tmp[622]*kernel[3]+tmp[623]*kernel[4]+tmp[624]*kernel[5]+tmp[722]*kernel[6]+tmp[723]*kernel[7]+tmp[724]*kernel[8];
				ans[624]<=tmp[523]*kernel[0]+tmp[524]*kernel[1]+tmp[525]*kernel[2]+tmp[623]*kernel[3]+tmp[624]*kernel[4]+tmp[625]*kernel[5]+tmp[723]*kernel[6]+tmp[724]*kernel[7]+tmp[725]*kernel[8];
				ans[625]<=tmp[524]*kernel[0]+tmp[525]*kernel[1]+tmp[526]*kernel[2]+tmp[624]*kernel[3]+tmp[625]*kernel[4]+tmp[626]*kernel[5]+tmp[724]*kernel[6]+tmp[725]*kernel[7]+tmp[726]*kernel[8];
				ans[626]<=tmp[525]*kernel[0]+tmp[526]*kernel[1]+tmp[527]*kernel[2]+tmp[625]*kernel[3]+tmp[626]*kernel[4]+tmp[627]*kernel[5]+tmp[725]*kernel[6]+tmp[726]*kernel[7]+tmp[727]*kernel[8];
				ans[627]<=tmp[526]*kernel[0]+tmp[527]*kernel[1]+tmp[528]*kernel[2]+tmp[626]*kernel[3]+tmp[627]*kernel[4]+tmp[628]*kernel[5]+tmp[726]*kernel[6]+tmp[727]*kernel[7]+tmp[728]*kernel[8];
				ans[628]<=tmp[527]*kernel[0]+tmp[528]*kernel[1]+tmp[529]*kernel[2]+tmp[627]*kernel[3]+tmp[628]*kernel[4]+tmp[629]*kernel[5]+tmp[727]*kernel[6]+tmp[728]*kernel[7]+tmp[729]*kernel[8];
				ans[629]<=tmp[528]*kernel[0]+tmp[529]*kernel[1]+tmp[530]*kernel[2]+tmp[628]*kernel[3]+tmp[629]*kernel[4]+tmp[630]*kernel[5]+tmp[728]*kernel[6]+tmp[729]*kernel[7]+tmp[730]*kernel[8];
				ans[630]<=tmp[529]*kernel[0]+tmp[530]*kernel[1]+tmp[531]*kernel[2]+tmp[629]*kernel[3]+tmp[630]*kernel[4]+tmp[631]*kernel[5]+tmp[729]*kernel[6]+tmp[730]*kernel[7]+tmp[731]*kernel[8];
				ans[631]<=tmp[530]*kernel[0]+tmp[531]*kernel[1]+tmp[532]*kernel[2]+tmp[630]*kernel[3]+tmp[631]*kernel[4]+tmp[632]*kernel[5]+tmp[730]*kernel[6]+tmp[731]*kernel[7]+tmp[732]*kernel[8];
				ans[632]<=tmp[531]*kernel[0]+tmp[532]*kernel[1]+tmp[533]*kernel[2]+tmp[631]*kernel[3]+tmp[632]*kernel[4]+tmp[633]*kernel[5]+tmp[731]*kernel[6]+tmp[732]*kernel[7]+tmp[733]*kernel[8];
				ans[633]<=tmp[532]*kernel[0]+tmp[533]*kernel[1]+tmp[534]*kernel[2]+tmp[632]*kernel[3]+tmp[633]*kernel[4]+tmp[634]*kernel[5]+tmp[732]*kernel[6]+tmp[733]*kernel[7]+tmp[734]*kernel[8];
				ans[634]<=tmp[533]*kernel[0]+tmp[534]*kernel[1]+tmp[535]*kernel[2]+tmp[633]*kernel[3]+tmp[634]*kernel[4]+tmp[635]*kernel[5]+tmp[733]*kernel[6]+tmp[734]*kernel[7]+tmp[735]*kernel[8];
				ans[635]<=tmp[534]*kernel[0]+tmp[535]*kernel[1]+tmp[536]*kernel[2]+tmp[634]*kernel[3]+tmp[635]*kernel[4]+tmp[636]*kernel[5]+tmp[734]*kernel[6]+tmp[735]*kernel[7]+tmp[736]*kernel[8];
				ans[636]<=tmp[535]*kernel[0]+tmp[536]*kernel[1]+tmp[537]*kernel[2]+tmp[635]*kernel[3]+tmp[636]*kernel[4]+tmp[637]*kernel[5]+tmp[735]*kernel[6]+tmp[736]*kernel[7]+tmp[737]*kernel[8];
				ans[637]<=tmp[536]*kernel[0]+tmp[537]*kernel[1]+tmp[538]*kernel[2]+tmp[636]*kernel[3]+tmp[637]*kernel[4]+tmp[638]*kernel[5]+tmp[736]*kernel[6]+tmp[737]*kernel[7]+tmp[738]*kernel[8];
				ans[638]<=tmp[537]*kernel[0]+tmp[538]*kernel[1]+tmp[539]*kernel[2]+tmp[637]*kernel[3]+tmp[638]*kernel[4]+tmp[639]*kernel[5]+tmp[737]*kernel[6]+tmp[738]*kernel[7]+tmp[739]*kernel[8];
				ans[639]<=tmp[538]*kernel[0]+tmp[539]*kernel[1]+tmp[540]*kernel[2]+tmp[638]*kernel[3]+tmp[639]*kernel[4]+tmp[640]*kernel[5]+tmp[738]*kernel[6]+tmp[739]*kernel[7]+tmp[740]*kernel[8];
				ans[640]<=tmp[539]*kernel[0]+tmp[540]*kernel[1]+tmp[541]*kernel[2]+tmp[639]*kernel[3]+tmp[640]*kernel[4]+tmp[641]*kernel[5]+tmp[739]*kernel[6]+tmp[740]*kernel[7]+tmp[741]*kernel[8];
				ans[641]<=tmp[540]*kernel[0]+tmp[541]*kernel[1]+tmp[542]*kernel[2]+tmp[640]*kernel[3]+tmp[641]*kernel[4]+tmp[642]*kernel[5]+tmp[740]*kernel[6]+tmp[741]*kernel[7]+tmp[742]*kernel[8];
				ans[642]<=tmp[541]*kernel[0]+tmp[542]*kernel[1]+tmp[543]*kernel[2]+tmp[641]*kernel[3]+tmp[642]*kernel[4]+tmp[643]*kernel[5]+tmp[741]*kernel[6]+tmp[742]*kernel[7]+tmp[743]*kernel[8];
				ans[643]<=tmp[542]*kernel[0]+tmp[543]*kernel[1]+tmp[544]*kernel[2]+tmp[642]*kernel[3]+tmp[643]*kernel[4]+tmp[644]*kernel[5]+tmp[742]*kernel[6]+tmp[743]*kernel[7]+tmp[744]*kernel[8];
				ans[644]<=tmp[543]*kernel[0]+tmp[544]*kernel[1]+tmp[545]*kernel[2]+tmp[643]*kernel[3]+tmp[644]*kernel[4]+tmp[645]*kernel[5]+tmp[743]*kernel[6]+tmp[744]*kernel[7]+tmp[745]*kernel[8];
				ans[645]<=tmp[544]*kernel[0]+tmp[545]*kernel[1]+tmp[546]*kernel[2]+tmp[644]*kernel[3]+tmp[645]*kernel[4]+tmp[646]*kernel[5]+tmp[744]*kernel[6]+tmp[745]*kernel[7]+tmp[746]*kernel[8];
				ans[646]<=tmp[545]*kernel[0]+tmp[546]*kernel[1]+tmp[547]*kernel[2]+tmp[645]*kernel[3]+tmp[646]*kernel[4]+tmp[647]*kernel[5]+tmp[745]*kernel[6]+tmp[746]*kernel[7]+tmp[747]*kernel[8];
				ans[647]<=tmp[546]*kernel[0]+tmp[547]*kernel[1]+tmp[548]*kernel[2]+tmp[646]*kernel[3]+tmp[647]*kernel[4]+tmp[648]*kernel[5]+tmp[746]*kernel[6]+tmp[747]*kernel[7]+tmp[748]*kernel[8];
				ans[648]<=tmp[547]*kernel[0]+tmp[548]*kernel[1]+tmp[549]*kernel[2]+tmp[647]*kernel[3]+tmp[648]*kernel[4]+tmp[649]*kernel[5]+tmp[747]*kernel[6]+tmp[748]*kernel[7]+tmp[749]*kernel[8];
				ans[649]<=tmp[548]*kernel[0]+tmp[549]*kernel[1]+tmp[550]*kernel[2]+tmp[648]*kernel[3]+tmp[649]*kernel[4]+tmp[650]*kernel[5]+tmp[748]*kernel[6]+tmp[749]*kernel[7]+tmp[750]*kernel[8];
				ans[650]<=tmp[549]*kernel[0]+tmp[550]*kernel[1]+tmp[551]*kernel[2]+tmp[649]*kernel[3]+tmp[650]*kernel[4]+tmp[651]*kernel[5]+tmp[749]*kernel[6]+tmp[750]*kernel[7]+tmp[751]*kernel[8];
				ans[651]<=tmp[550]*kernel[0]+tmp[551]*kernel[1]+tmp[552]*kernel[2]+tmp[650]*kernel[3]+tmp[651]*kernel[4]+tmp[652]*kernel[5]+tmp[750]*kernel[6]+tmp[751]*kernel[7]+tmp[752]*kernel[8];
				ans[652]<=tmp[551]*kernel[0]+tmp[552]*kernel[1]+tmp[553]*kernel[2]+tmp[651]*kernel[3]+tmp[652]*kernel[4]+tmp[653]*kernel[5]+tmp[751]*kernel[6]+tmp[752]*kernel[7]+tmp[753]*kernel[8];
				ans[653]<=tmp[552]*kernel[0]+tmp[553]*kernel[1]+tmp[554]*kernel[2]+tmp[652]*kernel[3]+tmp[653]*kernel[4]+tmp[654]*kernel[5]+tmp[752]*kernel[6]+tmp[753]*kernel[7]+tmp[754]*kernel[8];
				ans[654]<=tmp[553]*kernel[0]+tmp[554]*kernel[1]+tmp[555]*kernel[2]+tmp[653]*kernel[3]+tmp[654]*kernel[4]+tmp[655]*kernel[5]+tmp[753]*kernel[6]+tmp[754]*kernel[7]+tmp[755]*kernel[8];
				ans[655]<=tmp[554]*kernel[0]+tmp[555]*kernel[1]+tmp[556]*kernel[2]+tmp[654]*kernel[3]+tmp[655]*kernel[4]+tmp[656]*kernel[5]+tmp[754]*kernel[6]+tmp[755]*kernel[7]+tmp[756]*kernel[8];
				ans[656]<=tmp[555]*kernel[0]+tmp[556]*kernel[1]+tmp[557]*kernel[2]+tmp[655]*kernel[3]+tmp[656]*kernel[4]+tmp[657]*kernel[5]+tmp[755]*kernel[6]+tmp[756]*kernel[7]+tmp[757]*kernel[8];
				ans[657]<=tmp[556]*kernel[0]+tmp[557]*kernel[1]+tmp[558]*kernel[2]+tmp[656]*kernel[3]+tmp[657]*kernel[4]+tmp[658]*kernel[5]+tmp[756]*kernel[6]+tmp[757]*kernel[7]+tmp[758]*kernel[8];
				ans[658]<=tmp[557]*kernel[0]+tmp[558]*kernel[1]+tmp[559]*kernel[2]+tmp[657]*kernel[3]+tmp[658]*kernel[4]+tmp[659]*kernel[5]+tmp[757]*kernel[6]+tmp[758]*kernel[7]+tmp[759]*kernel[8];
				ans[659]<=tmp[558]*kernel[0]+tmp[559]*kernel[1]+tmp[560]*kernel[2]+tmp[658]*kernel[3]+tmp[659]*kernel[4]+tmp[660]*kernel[5]+tmp[758]*kernel[6]+tmp[759]*kernel[7]+tmp[760]*kernel[8];
				ans[660]<=tmp[559]*kernel[0]+tmp[560]*kernel[1]+tmp[561]*kernel[2]+tmp[659]*kernel[3]+tmp[660]*kernel[4]+tmp[661]*kernel[5]+tmp[759]*kernel[6]+tmp[760]*kernel[7]+tmp[761]*kernel[8];
				ans[661]<=tmp[560]*kernel[0]+tmp[561]*kernel[1]+tmp[562]*kernel[2]+tmp[660]*kernel[3]+tmp[661]*kernel[4]+tmp[662]*kernel[5]+tmp[760]*kernel[6]+tmp[761]*kernel[7]+tmp[762]*kernel[8];
				ans[662]<=tmp[561]*kernel[0]+tmp[562]*kernel[1]+tmp[563]*kernel[2]+tmp[661]*kernel[3]+tmp[662]*kernel[4]+tmp[663]*kernel[5]+tmp[761]*kernel[6]+tmp[762]*kernel[7]+tmp[763]*kernel[8];
				ans[663]<=tmp[562]*kernel[0]+tmp[563]*kernel[1]+tmp[564]*kernel[2]+tmp[662]*kernel[3]+tmp[663]*kernel[4]+tmp[664]*kernel[5]+tmp[762]*kernel[6]+tmp[763]*kernel[7]+tmp[764]*kernel[8];
				ans[664]<=tmp[563]*kernel[0]+tmp[564]*kernel[1]+tmp[565]*kernel[2]+tmp[663]*kernel[3]+tmp[664]*kernel[4]+tmp[665]*kernel[5]+tmp[763]*kernel[6]+tmp[764]*kernel[7]+tmp[765]*kernel[8];
				ans[665]<=tmp[564]*kernel[0]+tmp[565]*kernel[1]+tmp[566]*kernel[2]+tmp[664]*kernel[3]+tmp[665]*kernel[4]+tmp[666]*kernel[5]+tmp[764]*kernel[6]+tmp[765]*kernel[7]+tmp[766]*kernel[8];
				ans[666]<=tmp[565]*kernel[0]+tmp[566]*kernel[1]+tmp[567]*kernel[2]+tmp[665]*kernel[3]+tmp[666]*kernel[4]+tmp[667]*kernel[5]+tmp[765]*kernel[6]+tmp[766]*kernel[7]+tmp[767]*kernel[8];
				ans[667]<=tmp[566]*kernel[0]+tmp[567]*kernel[1]+tmp[568]*kernel[2]+tmp[666]*kernel[3]+tmp[667]*kernel[4]+tmp[668]*kernel[5]+tmp[766]*kernel[6]+tmp[767]*kernel[7]+tmp[768]*kernel[8];
				ans[668]<=tmp[567]*kernel[0]+tmp[568]*kernel[1]+tmp[569]*kernel[2]+tmp[667]*kernel[3]+tmp[668]*kernel[4]+tmp[669]*kernel[5]+tmp[767]*kernel[6]+tmp[768]*kernel[7]+tmp[769]*kernel[8];
				ans[669]<=tmp[568]*kernel[0]+tmp[569]*kernel[1]+tmp[570]*kernel[2]+tmp[668]*kernel[3]+tmp[669]*kernel[4]+tmp[670]*kernel[5]+tmp[768]*kernel[6]+tmp[769]*kernel[7]+tmp[770]*kernel[8];
				ans[670]<=tmp[569]*kernel[0]+tmp[570]*kernel[1]+tmp[571]*kernel[2]+tmp[669]*kernel[3]+tmp[670]*kernel[4]+tmp[671]*kernel[5]+tmp[769]*kernel[6]+tmp[770]*kernel[7]+tmp[771]*kernel[8];
				ans[671]<=tmp[570]*kernel[0]+tmp[571]*kernel[1]+tmp[572]*kernel[2]+tmp[670]*kernel[3]+tmp[671]*kernel[4]+tmp[672]*kernel[5]+tmp[770]*kernel[6]+tmp[771]*kernel[7]+tmp[772]*kernel[8];
				ans[672]<=tmp[571]*kernel[0]+tmp[572]*kernel[1]+tmp[573]*kernel[2]+tmp[671]*kernel[3]+tmp[672]*kernel[4]+tmp[673]*kernel[5]+tmp[771]*kernel[6]+tmp[772]*kernel[7]+tmp[773]*kernel[8];
				ans[673]<=tmp[572]*kernel[0]+tmp[573]*kernel[1]+tmp[574]*kernel[2]+tmp[672]*kernel[3]+tmp[673]*kernel[4]+tmp[674]*kernel[5]+tmp[772]*kernel[6]+tmp[773]*kernel[7]+tmp[774]*kernel[8];
				ans[674]<=tmp[573]*kernel[0]+tmp[574]*kernel[1]+tmp[575]*kernel[2]+tmp[673]*kernel[3]+tmp[674]*kernel[4]+tmp[675]*kernel[5]+tmp[773]*kernel[6]+tmp[774]*kernel[7]+tmp[775]*kernel[8];
				ans[675]<=tmp[574]*kernel[0]+tmp[575]*kernel[1]+tmp[576]*kernel[2]+tmp[674]*kernel[3]+tmp[675]*kernel[4]+tmp[676]*kernel[5]+tmp[774]*kernel[6]+tmp[775]*kernel[7]+tmp[776]*kernel[8];
				ans[676]<=tmp[575]*kernel[0]+tmp[576]*kernel[1]+tmp[577]*kernel[2]+tmp[675]*kernel[3]+tmp[676]*kernel[4]+tmp[677]*kernel[5]+tmp[775]*kernel[6]+tmp[776]*kernel[7]+tmp[777]*kernel[8];
				ans[677]<=tmp[576]*kernel[0]+tmp[577]*kernel[1]+tmp[578]*kernel[2]+tmp[676]*kernel[3]+tmp[677]*kernel[4]+tmp[678]*kernel[5]+tmp[776]*kernel[6]+tmp[777]*kernel[7]+tmp[778]*kernel[8];
				ans[678]<=tmp[577]*kernel[0]+tmp[578]*kernel[1]+tmp[579]*kernel[2]+tmp[677]*kernel[3]+tmp[678]*kernel[4]+tmp[679]*kernel[5]+tmp[777]*kernel[6]+tmp[778]*kernel[7]+tmp[779]*kernel[8];
				ans[679]<=tmp[578]*kernel[0]+tmp[579]*kernel[1]+tmp[580]*kernel[2]+tmp[678]*kernel[3]+tmp[679]*kernel[4]+tmp[680]*kernel[5]+tmp[778]*kernel[6]+tmp[779]*kernel[7]+tmp[780]*kernel[8];
				ans[680]<=tmp[579]*kernel[0]+tmp[580]*kernel[1]+tmp[581]*kernel[2]+tmp[679]*kernel[3]+tmp[680]*kernel[4]+tmp[681]*kernel[5]+tmp[779]*kernel[6]+tmp[780]*kernel[7]+tmp[781]*kernel[8];
				ans[681]<=tmp[580]*kernel[0]+tmp[581]*kernel[1]+tmp[582]*kernel[2]+tmp[680]*kernel[3]+tmp[681]*kernel[4]+tmp[682]*kernel[5]+tmp[780]*kernel[6]+tmp[781]*kernel[7]+tmp[782]*kernel[8];
				ans[682]<=tmp[581]*kernel[0]+tmp[582]*kernel[1]+tmp[583]*kernel[2]+tmp[681]*kernel[3]+tmp[682]*kernel[4]+tmp[683]*kernel[5]+tmp[781]*kernel[6]+tmp[782]*kernel[7]+tmp[783]*kernel[8];
				ans[683]<=tmp[582]*kernel[0]+tmp[583]*kernel[1]+tmp[584]*kernel[2]+tmp[682]*kernel[3]+tmp[683]*kernel[4]+tmp[684]*kernel[5]+tmp[782]*kernel[6]+tmp[783]*kernel[7]+tmp[784]*kernel[8];
				ans[684]<=tmp[583]*kernel[0]+tmp[584]*kernel[1]+tmp[585]*kernel[2]+tmp[683]*kernel[3]+tmp[684]*kernel[4]+tmp[685]*kernel[5]+tmp[783]*kernel[6]+tmp[784]*kernel[7]+tmp[785]*kernel[8];
				ans[685]<=tmp[584]*kernel[0]+tmp[585]*kernel[1]+tmp[586]*kernel[2]+tmp[684]*kernel[3]+tmp[685]*kernel[4]+tmp[686]*kernel[5]+tmp[784]*kernel[6]+tmp[785]*kernel[7]+tmp[786]*kernel[8];
				ans[686]<=tmp[585]*kernel[0]+tmp[586]*kernel[1]+tmp[587]*kernel[2]+tmp[685]*kernel[3]+tmp[686]*kernel[4]+tmp[687]*kernel[5]+tmp[785]*kernel[6]+tmp[786]*kernel[7]+tmp[787]*kernel[8];
				ans[687]<=tmp[586]*kernel[0]+tmp[587]*kernel[1]+tmp[588]*kernel[2]+tmp[686]*kernel[3]+tmp[687]*kernel[4]+tmp[688]*kernel[5]+tmp[786]*kernel[6]+tmp[787]*kernel[7]+tmp[788]*kernel[8];
				ans[688]<=tmp[587]*kernel[0]+tmp[588]*kernel[1]+tmp[589]*kernel[2]+tmp[687]*kernel[3]+tmp[688]*kernel[4]+tmp[689]*kernel[5]+tmp[787]*kernel[6]+tmp[788]*kernel[7]+tmp[789]*kernel[8];
				ans[689]<=tmp[588]*kernel[0]+tmp[589]*kernel[1]+tmp[590]*kernel[2]+tmp[688]*kernel[3]+tmp[689]*kernel[4]+tmp[690]*kernel[5]+tmp[788]*kernel[6]+tmp[789]*kernel[7]+tmp[790]*kernel[8];
				ans[690]<=tmp[589]*kernel[0]+tmp[590]*kernel[1]+tmp[591]*kernel[2]+tmp[689]*kernel[3]+tmp[690]*kernel[4]+tmp[691]*kernel[5]+tmp[789]*kernel[6]+tmp[790]*kernel[7]+tmp[791]*kernel[8];
				ans[691]<=tmp[590]*kernel[0]+tmp[591]*kernel[1]+tmp[592]*kernel[2]+tmp[690]*kernel[3]+tmp[691]*kernel[4]+tmp[692]*kernel[5]+tmp[790]*kernel[6]+tmp[791]*kernel[7]+tmp[792]*kernel[8];
				ans[692]<=tmp[591]*kernel[0]+tmp[592]*kernel[1]+tmp[593]*kernel[2]+tmp[691]*kernel[3]+tmp[692]*kernel[4]+tmp[693]*kernel[5]+tmp[791]*kernel[6]+tmp[792]*kernel[7]+tmp[793]*kernel[8];
				ans[693]<=tmp[592]*kernel[0]+tmp[593]*kernel[1]+tmp[594]*kernel[2]+tmp[692]*kernel[3]+tmp[693]*kernel[4]+tmp[694]*kernel[5]+tmp[792]*kernel[6]+tmp[793]*kernel[7]+tmp[794]*kernel[8];
				ans[694]<=tmp[593]*kernel[0]+tmp[594]*kernel[1]+tmp[595]*kernel[2]+tmp[693]*kernel[3]+tmp[694]*kernel[4]+tmp[695]*kernel[5]+tmp[793]*kernel[6]+tmp[794]*kernel[7]+tmp[795]*kernel[8];
				ans[695]<=tmp[594]*kernel[0]+tmp[595]*kernel[1]+tmp[596]*kernel[2]+tmp[694]*kernel[3]+tmp[695]*kernel[4]+tmp[696]*kernel[5]+tmp[794]*kernel[6]+tmp[795]*kernel[7]+tmp[796]*kernel[8];
				ans[696]<=tmp[595]*kernel[0]+tmp[596]*kernel[1]+tmp[597]*kernel[2]+tmp[695]*kernel[3]+tmp[696]*kernel[4]+tmp[697]*kernel[5]+tmp[795]*kernel[6]+tmp[796]*kernel[7]+tmp[797]*kernel[8];
				ans[697]<=tmp[596]*kernel[0]+tmp[597]*kernel[1]+tmp[598]*kernel[2]+tmp[696]*kernel[3]+tmp[697]*kernel[4]+tmp[698]*kernel[5]+tmp[796]*kernel[6]+tmp[797]*kernel[7]+tmp[798]*kernel[8];
				ans[698]<=tmp[597]*kernel[0]+tmp[598]*kernel[1]+tmp[599]*kernel[2]+tmp[697]*kernel[3]+tmp[698]*kernel[4]+tmp[699]*kernel[5]+tmp[797]*kernel[6]+tmp[798]*kernel[7]+tmp[799]*kernel[8];
				ans[699]<=tmp[598]*kernel[0]+tmp[599]*kernel[1]+tmp[698]*kernel[3]+tmp[699]*kernel[4]+tmp[798]*kernel[6]+tmp[799]*kernel[7];
				ans[700]<=tmp[600]*kernel[1]+tmp[601]*kernel[2]+tmp[700]*kernel[4]+tmp[701]*kernel[5]+tmp[800]*kernel[7]+tmp[801]*kernel[8];
				ans[701]<=tmp[600]*kernel[0]+tmp[601]*kernel[1]+tmp[602]*kernel[2]+tmp[700]*kernel[3]+tmp[701]*kernel[4]+tmp[702]*kernel[5]+tmp[800]*kernel[6]+tmp[801]*kernel[7]+tmp[802]*kernel[8];
				ans[702]<=tmp[601]*kernel[0]+tmp[602]*kernel[1]+tmp[603]*kernel[2]+tmp[701]*kernel[3]+tmp[702]*kernel[4]+tmp[703]*kernel[5]+tmp[801]*kernel[6]+tmp[802]*kernel[7]+tmp[803]*kernel[8];
				ans[703]<=tmp[602]*kernel[0]+tmp[603]*kernel[1]+tmp[604]*kernel[2]+tmp[702]*kernel[3]+tmp[703]*kernel[4]+tmp[704]*kernel[5]+tmp[802]*kernel[6]+tmp[803]*kernel[7]+tmp[804]*kernel[8];
				ans[704]<=tmp[603]*kernel[0]+tmp[604]*kernel[1]+tmp[605]*kernel[2]+tmp[703]*kernel[3]+tmp[704]*kernel[4]+tmp[705]*kernel[5]+tmp[803]*kernel[6]+tmp[804]*kernel[7]+tmp[805]*kernel[8];
				ans[705]<=tmp[604]*kernel[0]+tmp[605]*kernel[1]+tmp[606]*kernel[2]+tmp[704]*kernel[3]+tmp[705]*kernel[4]+tmp[706]*kernel[5]+tmp[804]*kernel[6]+tmp[805]*kernel[7]+tmp[806]*kernel[8];
				ans[706]<=tmp[605]*kernel[0]+tmp[606]*kernel[1]+tmp[607]*kernel[2]+tmp[705]*kernel[3]+tmp[706]*kernel[4]+tmp[707]*kernel[5]+tmp[805]*kernel[6]+tmp[806]*kernel[7]+tmp[807]*kernel[8];
				ans[707]<=tmp[606]*kernel[0]+tmp[607]*kernel[1]+tmp[608]*kernel[2]+tmp[706]*kernel[3]+tmp[707]*kernel[4]+tmp[708]*kernel[5]+tmp[806]*kernel[6]+tmp[807]*kernel[7]+tmp[808]*kernel[8];
				ans[708]<=tmp[607]*kernel[0]+tmp[608]*kernel[1]+tmp[609]*kernel[2]+tmp[707]*kernel[3]+tmp[708]*kernel[4]+tmp[709]*kernel[5]+tmp[807]*kernel[6]+tmp[808]*kernel[7]+tmp[809]*kernel[8];
				ans[709]<=tmp[608]*kernel[0]+tmp[609]*kernel[1]+tmp[610]*kernel[2]+tmp[708]*kernel[3]+tmp[709]*kernel[4]+tmp[710]*kernel[5]+tmp[808]*kernel[6]+tmp[809]*kernel[7]+tmp[810]*kernel[8];
				ans[710]<=tmp[609]*kernel[0]+tmp[610]*kernel[1]+tmp[611]*kernel[2]+tmp[709]*kernel[3]+tmp[710]*kernel[4]+tmp[711]*kernel[5]+tmp[809]*kernel[6]+tmp[810]*kernel[7]+tmp[811]*kernel[8];
				ans[711]<=tmp[610]*kernel[0]+tmp[611]*kernel[1]+tmp[612]*kernel[2]+tmp[710]*kernel[3]+tmp[711]*kernel[4]+tmp[712]*kernel[5]+tmp[810]*kernel[6]+tmp[811]*kernel[7]+tmp[812]*kernel[8];
				ans[712]<=tmp[611]*kernel[0]+tmp[612]*kernel[1]+tmp[613]*kernel[2]+tmp[711]*kernel[3]+tmp[712]*kernel[4]+tmp[713]*kernel[5]+tmp[811]*kernel[6]+tmp[812]*kernel[7]+tmp[813]*kernel[8];
				ans[713]<=tmp[612]*kernel[0]+tmp[613]*kernel[1]+tmp[614]*kernel[2]+tmp[712]*kernel[3]+tmp[713]*kernel[4]+tmp[714]*kernel[5]+tmp[812]*kernel[6]+tmp[813]*kernel[7]+tmp[814]*kernel[8];
				ans[714]<=tmp[613]*kernel[0]+tmp[614]*kernel[1]+tmp[615]*kernel[2]+tmp[713]*kernel[3]+tmp[714]*kernel[4]+tmp[715]*kernel[5]+tmp[813]*kernel[6]+tmp[814]*kernel[7]+tmp[815]*kernel[8];
				ans[715]<=tmp[614]*kernel[0]+tmp[615]*kernel[1]+tmp[616]*kernel[2]+tmp[714]*kernel[3]+tmp[715]*kernel[4]+tmp[716]*kernel[5]+tmp[814]*kernel[6]+tmp[815]*kernel[7]+tmp[816]*kernel[8];
				ans[716]<=tmp[615]*kernel[0]+tmp[616]*kernel[1]+tmp[617]*kernel[2]+tmp[715]*kernel[3]+tmp[716]*kernel[4]+tmp[717]*kernel[5]+tmp[815]*kernel[6]+tmp[816]*kernel[7]+tmp[817]*kernel[8];
				ans[717]<=tmp[616]*kernel[0]+tmp[617]*kernel[1]+tmp[618]*kernel[2]+tmp[716]*kernel[3]+tmp[717]*kernel[4]+tmp[718]*kernel[5]+tmp[816]*kernel[6]+tmp[817]*kernel[7]+tmp[818]*kernel[8];
				ans[718]<=tmp[617]*kernel[0]+tmp[618]*kernel[1]+tmp[619]*kernel[2]+tmp[717]*kernel[3]+tmp[718]*kernel[4]+tmp[719]*kernel[5]+tmp[817]*kernel[6]+tmp[818]*kernel[7]+tmp[819]*kernel[8];
				ans[719]<=tmp[618]*kernel[0]+tmp[619]*kernel[1]+tmp[620]*kernel[2]+tmp[718]*kernel[3]+tmp[719]*kernel[4]+tmp[720]*kernel[5]+tmp[818]*kernel[6]+tmp[819]*kernel[7]+tmp[820]*kernel[8];
				ans[720]<=tmp[619]*kernel[0]+tmp[620]*kernel[1]+tmp[621]*kernel[2]+tmp[719]*kernel[3]+tmp[720]*kernel[4]+tmp[721]*kernel[5]+tmp[819]*kernel[6]+tmp[820]*kernel[7]+tmp[821]*kernel[8];
				ans[721]<=tmp[620]*kernel[0]+tmp[621]*kernel[1]+tmp[622]*kernel[2]+tmp[720]*kernel[3]+tmp[721]*kernel[4]+tmp[722]*kernel[5]+tmp[820]*kernel[6]+tmp[821]*kernel[7]+tmp[822]*kernel[8];
				ans[722]<=tmp[621]*kernel[0]+tmp[622]*kernel[1]+tmp[623]*kernel[2]+tmp[721]*kernel[3]+tmp[722]*kernel[4]+tmp[723]*kernel[5]+tmp[821]*kernel[6]+tmp[822]*kernel[7]+tmp[823]*kernel[8];
				ans[723]<=tmp[622]*kernel[0]+tmp[623]*kernel[1]+tmp[624]*kernel[2]+tmp[722]*kernel[3]+tmp[723]*kernel[4]+tmp[724]*kernel[5]+tmp[822]*kernel[6]+tmp[823]*kernel[7]+tmp[824]*kernel[8];
				ans[724]<=tmp[623]*kernel[0]+tmp[624]*kernel[1]+tmp[625]*kernel[2]+tmp[723]*kernel[3]+tmp[724]*kernel[4]+tmp[725]*kernel[5]+tmp[823]*kernel[6]+tmp[824]*kernel[7]+tmp[825]*kernel[8];
				ans[725]<=tmp[624]*kernel[0]+tmp[625]*kernel[1]+tmp[626]*kernel[2]+tmp[724]*kernel[3]+tmp[725]*kernel[4]+tmp[726]*kernel[5]+tmp[824]*kernel[6]+tmp[825]*kernel[7]+tmp[826]*kernel[8];
				ans[726]<=tmp[625]*kernel[0]+tmp[626]*kernel[1]+tmp[627]*kernel[2]+tmp[725]*kernel[3]+tmp[726]*kernel[4]+tmp[727]*kernel[5]+tmp[825]*kernel[6]+tmp[826]*kernel[7]+tmp[827]*kernel[8];
				ans[727]<=tmp[626]*kernel[0]+tmp[627]*kernel[1]+tmp[628]*kernel[2]+tmp[726]*kernel[3]+tmp[727]*kernel[4]+tmp[728]*kernel[5]+tmp[826]*kernel[6]+tmp[827]*kernel[7]+tmp[828]*kernel[8];
				ans[728]<=tmp[627]*kernel[0]+tmp[628]*kernel[1]+tmp[629]*kernel[2]+tmp[727]*kernel[3]+tmp[728]*kernel[4]+tmp[729]*kernel[5]+tmp[827]*kernel[6]+tmp[828]*kernel[7]+tmp[829]*kernel[8];
				ans[729]<=tmp[628]*kernel[0]+tmp[629]*kernel[1]+tmp[630]*kernel[2]+tmp[728]*kernel[3]+tmp[729]*kernel[4]+tmp[730]*kernel[5]+tmp[828]*kernel[6]+tmp[829]*kernel[7]+tmp[830]*kernel[8];
				ans[730]<=tmp[629]*kernel[0]+tmp[630]*kernel[1]+tmp[631]*kernel[2]+tmp[729]*kernel[3]+tmp[730]*kernel[4]+tmp[731]*kernel[5]+tmp[829]*kernel[6]+tmp[830]*kernel[7]+tmp[831]*kernel[8];
				ans[731]<=tmp[630]*kernel[0]+tmp[631]*kernel[1]+tmp[632]*kernel[2]+tmp[730]*kernel[3]+tmp[731]*kernel[4]+tmp[732]*kernel[5]+tmp[830]*kernel[6]+tmp[831]*kernel[7]+tmp[832]*kernel[8];
				ans[732]<=tmp[631]*kernel[0]+tmp[632]*kernel[1]+tmp[633]*kernel[2]+tmp[731]*kernel[3]+tmp[732]*kernel[4]+tmp[733]*kernel[5]+tmp[831]*kernel[6]+tmp[832]*kernel[7]+tmp[833]*kernel[8];
				ans[733]<=tmp[632]*kernel[0]+tmp[633]*kernel[1]+tmp[634]*kernel[2]+tmp[732]*kernel[3]+tmp[733]*kernel[4]+tmp[734]*kernel[5]+tmp[832]*kernel[6]+tmp[833]*kernel[7]+tmp[834]*kernel[8];
				ans[734]<=tmp[633]*kernel[0]+tmp[634]*kernel[1]+tmp[635]*kernel[2]+tmp[733]*kernel[3]+tmp[734]*kernel[4]+tmp[735]*kernel[5]+tmp[833]*kernel[6]+tmp[834]*kernel[7]+tmp[835]*kernel[8];
				ans[735]<=tmp[634]*kernel[0]+tmp[635]*kernel[1]+tmp[636]*kernel[2]+tmp[734]*kernel[3]+tmp[735]*kernel[4]+tmp[736]*kernel[5]+tmp[834]*kernel[6]+tmp[835]*kernel[7]+tmp[836]*kernel[8];
				ans[736]<=tmp[635]*kernel[0]+tmp[636]*kernel[1]+tmp[637]*kernel[2]+tmp[735]*kernel[3]+tmp[736]*kernel[4]+tmp[737]*kernel[5]+tmp[835]*kernel[6]+tmp[836]*kernel[7]+tmp[837]*kernel[8];
				ans[737]<=tmp[636]*kernel[0]+tmp[637]*kernel[1]+tmp[638]*kernel[2]+tmp[736]*kernel[3]+tmp[737]*kernel[4]+tmp[738]*kernel[5]+tmp[836]*kernel[6]+tmp[837]*kernel[7]+tmp[838]*kernel[8];
				ans[738]<=tmp[637]*kernel[0]+tmp[638]*kernel[1]+tmp[639]*kernel[2]+tmp[737]*kernel[3]+tmp[738]*kernel[4]+tmp[739]*kernel[5]+tmp[837]*kernel[6]+tmp[838]*kernel[7]+tmp[839]*kernel[8];
				ans[739]<=tmp[638]*kernel[0]+tmp[639]*kernel[1]+tmp[640]*kernel[2]+tmp[738]*kernel[3]+tmp[739]*kernel[4]+tmp[740]*kernel[5]+tmp[838]*kernel[6]+tmp[839]*kernel[7]+tmp[840]*kernel[8];
				ans[740]<=tmp[639]*kernel[0]+tmp[640]*kernel[1]+tmp[641]*kernel[2]+tmp[739]*kernel[3]+tmp[740]*kernel[4]+tmp[741]*kernel[5]+tmp[839]*kernel[6]+tmp[840]*kernel[7]+tmp[841]*kernel[8];
				ans[741]<=tmp[640]*kernel[0]+tmp[641]*kernel[1]+tmp[642]*kernel[2]+tmp[740]*kernel[3]+tmp[741]*kernel[4]+tmp[742]*kernel[5]+tmp[840]*kernel[6]+tmp[841]*kernel[7]+tmp[842]*kernel[8];
				ans[742]<=tmp[641]*kernel[0]+tmp[642]*kernel[1]+tmp[643]*kernel[2]+tmp[741]*kernel[3]+tmp[742]*kernel[4]+tmp[743]*kernel[5]+tmp[841]*kernel[6]+tmp[842]*kernel[7]+tmp[843]*kernel[8];
				ans[743]<=tmp[642]*kernel[0]+tmp[643]*kernel[1]+tmp[644]*kernel[2]+tmp[742]*kernel[3]+tmp[743]*kernel[4]+tmp[744]*kernel[5]+tmp[842]*kernel[6]+tmp[843]*kernel[7]+tmp[844]*kernel[8];
				ans[744]<=tmp[643]*kernel[0]+tmp[644]*kernel[1]+tmp[645]*kernel[2]+tmp[743]*kernel[3]+tmp[744]*kernel[4]+tmp[745]*kernel[5]+tmp[843]*kernel[6]+tmp[844]*kernel[7]+tmp[845]*kernel[8];
				ans[745]<=tmp[644]*kernel[0]+tmp[645]*kernel[1]+tmp[646]*kernel[2]+tmp[744]*kernel[3]+tmp[745]*kernel[4]+tmp[746]*kernel[5]+tmp[844]*kernel[6]+tmp[845]*kernel[7]+tmp[846]*kernel[8];
				ans[746]<=tmp[645]*kernel[0]+tmp[646]*kernel[1]+tmp[647]*kernel[2]+tmp[745]*kernel[3]+tmp[746]*kernel[4]+tmp[747]*kernel[5]+tmp[845]*kernel[6]+tmp[846]*kernel[7]+tmp[847]*kernel[8];
				ans[747]<=tmp[646]*kernel[0]+tmp[647]*kernel[1]+tmp[648]*kernel[2]+tmp[746]*kernel[3]+tmp[747]*kernel[4]+tmp[748]*kernel[5]+tmp[846]*kernel[6]+tmp[847]*kernel[7]+tmp[848]*kernel[8];
				ans[748]<=tmp[647]*kernel[0]+tmp[648]*kernel[1]+tmp[649]*kernel[2]+tmp[747]*kernel[3]+tmp[748]*kernel[4]+tmp[749]*kernel[5]+tmp[847]*kernel[6]+tmp[848]*kernel[7]+tmp[849]*kernel[8];
				ans[749]<=tmp[648]*kernel[0]+tmp[649]*kernel[1]+tmp[650]*kernel[2]+tmp[748]*kernel[3]+tmp[749]*kernel[4]+tmp[750]*kernel[5]+tmp[848]*kernel[6]+tmp[849]*kernel[7]+tmp[850]*kernel[8];
				ans[750]<=tmp[649]*kernel[0]+tmp[650]*kernel[1]+tmp[651]*kernel[2]+tmp[749]*kernel[3]+tmp[750]*kernel[4]+tmp[751]*kernel[5]+tmp[849]*kernel[6]+tmp[850]*kernel[7]+tmp[851]*kernel[8];
				ans[751]<=tmp[650]*kernel[0]+tmp[651]*kernel[1]+tmp[652]*kernel[2]+tmp[750]*kernel[3]+tmp[751]*kernel[4]+tmp[752]*kernel[5]+tmp[850]*kernel[6]+tmp[851]*kernel[7]+tmp[852]*kernel[8];
				ans[752]<=tmp[651]*kernel[0]+tmp[652]*kernel[1]+tmp[653]*kernel[2]+tmp[751]*kernel[3]+tmp[752]*kernel[4]+tmp[753]*kernel[5]+tmp[851]*kernel[6]+tmp[852]*kernel[7]+tmp[853]*kernel[8];
				ans[753]<=tmp[652]*kernel[0]+tmp[653]*kernel[1]+tmp[654]*kernel[2]+tmp[752]*kernel[3]+tmp[753]*kernel[4]+tmp[754]*kernel[5]+tmp[852]*kernel[6]+tmp[853]*kernel[7]+tmp[854]*kernel[8];
				ans[754]<=tmp[653]*kernel[0]+tmp[654]*kernel[1]+tmp[655]*kernel[2]+tmp[753]*kernel[3]+tmp[754]*kernel[4]+tmp[755]*kernel[5]+tmp[853]*kernel[6]+tmp[854]*kernel[7]+tmp[855]*kernel[8];
				ans[755]<=tmp[654]*kernel[0]+tmp[655]*kernel[1]+tmp[656]*kernel[2]+tmp[754]*kernel[3]+tmp[755]*kernel[4]+tmp[756]*kernel[5]+tmp[854]*kernel[6]+tmp[855]*kernel[7]+tmp[856]*kernel[8];
				ans[756]<=tmp[655]*kernel[0]+tmp[656]*kernel[1]+tmp[657]*kernel[2]+tmp[755]*kernel[3]+tmp[756]*kernel[4]+tmp[757]*kernel[5]+tmp[855]*kernel[6]+tmp[856]*kernel[7]+tmp[857]*kernel[8];
				ans[757]<=tmp[656]*kernel[0]+tmp[657]*kernel[1]+tmp[658]*kernel[2]+tmp[756]*kernel[3]+tmp[757]*kernel[4]+tmp[758]*kernel[5]+tmp[856]*kernel[6]+tmp[857]*kernel[7]+tmp[858]*kernel[8];
				ans[758]<=tmp[657]*kernel[0]+tmp[658]*kernel[1]+tmp[659]*kernel[2]+tmp[757]*kernel[3]+tmp[758]*kernel[4]+tmp[759]*kernel[5]+tmp[857]*kernel[6]+tmp[858]*kernel[7]+tmp[859]*kernel[8];
				ans[759]<=tmp[658]*kernel[0]+tmp[659]*kernel[1]+tmp[660]*kernel[2]+tmp[758]*kernel[3]+tmp[759]*kernel[4]+tmp[760]*kernel[5]+tmp[858]*kernel[6]+tmp[859]*kernel[7]+tmp[860]*kernel[8];
				ans[760]<=tmp[659]*kernel[0]+tmp[660]*kernel[1]+tmp[661]*kernel[2]+tmp[759]*kernel[3]+tmp[760]*kernel[4]+tmp[761]*kernel[5]+tmp[859]*kernel[6]+tmp[860]*kernel[7]+tmp[861]*kernel[8];
				ans[761]<=tmp[660]*kernel[0]+tmp[661]*kernel[1]+tmp[662]*kernel[2]+tmp[760]*kernel[3]+tmp[761]*kernel[4]+tmp[762]*kernel[5]+tmp[860]*kernel[6]+tmp[861]*kernel[7]+tmp[862]*kernel[8];
				ans[762]<=tmp[661]*kernel[0]+tmp[662]*kernel[1]+tmp[663]*kernel[2]+tmp[761]*kernel[3]+tmp[762]*kernel[4]+tmp[763]*kernel[5]+tmp[861]*kernel[6]+tmp[862]*kernel[7]+tmp[863]*kernel[8];
				ans[763]<=tmp[662]*kernel[0]+tmp[663]*kernel[1]+tmp[664]*kernel[2]+tmp[762]*kernel[3]+tmp[763]*kernel[4]+tmp[764]*kernel[5]+tmp[862]*kernel[6]+tmp[863]*kernel[7]+tmp[864]*kernel[8];
				ans[764]<=tmp[663]*kernel[0]+tmp[664]*kernel[1]+tmp[665]*kernel[2]+tmp[763]*kernel[3]+tmp[764]*kernel[4]+tmp[765]*kernel[5]+tmp[863]*kernel[6]+tmp[864]*kernel[7]+tmp[865]*kernel[8];
				ans[765]<=tmp[664]*kernel[0]+tmp[665]*kernel[1]+tmp[666]*kernel[2]+tmp[764]*kernel[3]+tmp[765]*kernel[4]+tmp[766]*kernel[5]+tmp[864]*kernel[6]+tmp[865]*kernel[7]+tmp[866]*kernel[8];
				ans[766]<=tmp[665]*kernel[0]+tmp[666]*kernel[1]+tmp[667]*kernel[2]+tmp[765]*kernel[3]+tmp[766]*kernel[4]+tmp[767]*kernel[5]+tmp[865]*kernel[6]+tmp[866]*kernel[7]+tmp[867]*kernel[8];
				ans[767]<=tmp[666]*kernel[0]+tmp[667]*kernel[1]+tmp[668]*kernel[2]+tmp[766]*kernel[3]+tmp[767]*kernel[4]+tmp[768]*kernel[5]+tmp[866]*kernel[6]+tmp[867]*kernel[7]+tmp[868]*kernel[8];
				ans[768]<=tmp[667]*kernel[0]+tmp[668]*kernel[1]+tmp[669]*kernel[2]+tmp[767]*kernel[3]+tmp[768]*kernel[4]+tmp[769]*kernel[5]+tmp[867]*kernel[6]+tmp[868]*kernel[7]+tmp[869]*kernel[8];
				ans[769]<=tmp[668]*kernel[0]+tmp[669]*kernel[1]+tmp[670]*kernel[2]+tmp[768]*kernel[3]+tmp[769]*kernel[4]+tmp[770]*kernel[5]+tmp[868]*kernel[6]+tmp[869]*kernel[7]+tmp[870]*kernel[8];
				ans[770]<=tmp[669]*kernel[0]+tmp[670]*kernel[1]+tmp[671]*kernel[2]+tmp[769]*kernel[3]+tmp[770]*kernel[4]+tmp[771]*kernel[5]+tmp[869]*kernel[6]+tmp[870]*kernel[7]+tmp[871]*kernel[8];
				ans[771]<=tmp[670]*kernel[0]+tmp[671]*kernel[1]+tmp[672]*kernel[2]+tmp[770]*kernel[3]+tmp[771]*kernel[4]+tmp[772]*kernel[5]+tmp[870]*kernel[6]+tmp[871]*kernel[7]+tmp[872]*kernel[8];
				ans[772]<=tmp[671]*kernel[0]+tmp[672]*kernel[1]+tmp[673]*kernel[2]+tmp[771]*kernel[3]+tmp[772]*kernel[4]+tmp[773]*kernel[5]+tmp[871]*kernel[6]+tmp[872]*kernel[7]+tmp[873]*kernel[8];
				ans[773]<=tmp[672]*kernel[0]+tmp[673]*kernel[1]+tmp[674]*kernel[2]+tmp[772]*kernel[3]+tmp[773]*kernel[4]+tmp[774]*kernel[5]+tmp[872]*kernel[6]+tmp[873]*kernel[7]+tmp[874]*kernel[8];
				ans[774]<=tmp[673]*kernel[0]+tmp[674]*kernel[1]+tmp[675]*kernel[2]+tmp[773]*kernel[3]+tmp[774]*kernel[4]+tmp[775]*kernel[5]+tmp[873]*kernel[6]+tmp[874]*kernel[7]+tmp[875]*kernel[8];
				ans[775]<=tmp[674]*kernel[0]+tmp[675]*kernel[1]+tmp[676]*kernel[2]+tmp[774]*kernel[3]+tmp[775]*kernel[4]+tmp[776]*kernel[5]+tmp[874]*kernel[6]+tmp[875]*kernel[7]+tmp[876]*kernel[8];
				ans[776]<=tmp[675]*kernel[0]+tmp[676]*kernel[1]+tmp[677]*kernel[2]+tmp[775]*kernel[3]+tmp[776]*kernel[4]+tmp[777]*kernel[5]+tmp[875]*kernel[6]+tmp[876]*kernel[7]+tmp[877]*kernel[8];
				ans[777]<=tmp[676]*kernel[0]+tmp[677]*kernel[1]+tmp[678]*kernel[2]+tmp[776]*kernel[3]+tmp[777]*kernel[4]+tmp[778]*kernel[5]+tmp[876]*kernel[6]+tmp[877]*kernel[7]+tmp[878]*kernel[8];
				ans[778]<=tmp[677]*kernel[0]+tmp[678]*kernel[1]+tmp[679]*kernel[2]+tmp[777]*kernel[3]+tmp[778]*kernel[4]+tmp[779]*kernel[5]+tmp[877]*kernel[6]+tmp[878]*kernel[7]+tmp[879]*kernel[8];
				ans[779]<=tmp[678]*kernel[0]+tmp[679]*kernel[1]+tmp[680]*kernel[2]+tmp[778]*kernel[3]+tmp[779]*kernel[4]+tmp[780]*kernel[5]+tmp[878]*kernel[6]+tmp[879]*kernel[7]+tmp[880]*kernel[8];
				ans[780]<=tmp[679]*kernel[0]+tmp[680]*kernel[1]+tmp[681]*kernel[2]+tmp[779]*kernel[3]+tmp[780]*kernel[4]+tmp[781]*kernel[5]+tmp[879]*kernel[6]+tmp[880]*kernel[7]+tmp[881]*kernel[8];
				ans[781]<=tmp[680]*kernel[0]+tmp[681]*kernel[1]+tmp[682]*kernel[2]+tmp[780]*kernel[3]+tmp[781]*kernel[4]+tmp[782]*kernel[5]+tmp[880]*kernel[6]+tmp[881]*kernel[7]+tmp[882]*kernel[8];
				ans[782]<=tmp[681]*kernel[0]+tmp[682]*kernel[1]+tmp[683]*kernel[2]+tmp[781]*kernel[3]+tmp[782]*kernel[4]+tmp[783]*kernel[5]+tmp[881]*kernel[6]+tmp[882]*kernel[7]+tmp[883]*kernel[8];
				ans[783]<=tmp[682]*kernel[0]+tmp[683]*kernel[1]+tmp[684]*kernel[2]+tmp[782]*kernel[3]+tmp[783]*kernel[4]+tmp[784]*kernel[5]+tmp[882]*kernel[6]+tmp[883]*kernel[7]+tmp[884]*kernel[8];
				ans[784]<=tmp[683]*kernel[0]+tmp[684]*kernel[1]+tmp[685]*kernel[2]+tmp[783]*kernel[3]+tmp[784]*kernel[4]+tmp[785]*kernel[5]+tmp[883]*kernel[6]+tmp[884]*kernel[7]+tmp[885]*kernel[8];
				ans[785]<=tmp[684]*kernel[0]+tmp[685]*kernel[1]+tmp[686]*kernel[2]+tmp[784]*kernel[3]+tmp[785]*kernel[4]+tmp[786]*kernel[5]+tmp[884]*kernel[6]+tmp[885]*kernel[7]+tmp[886]*kernel[8];
				ans[786]<=tmp[685]*kernel[0]+tmp[686]*kernel[1]+tmp[687]*kernel[2]+tmp[785]*kernel[3]+tmp[786]*kernel[4]+tmp[787]*kernel[5]+tmp[885]*kernel[6]+tmp[886]*kernel[7]+tmp[887]*kernel[8];
				ans[787]<=tmp[686]*kernel[0]+tmp[687]*kernel[1]+tmp[688]*kernel[2]+tmp[786]*kernel[3]+tmp[787]*kernel[4]+tmp[788]*kernel[5]+tmp[886]*kernel[6]+tmp[887]*kernel[7]+tmp[888]*kernel[8];
				ans[788]<=tmp[687]*kernel[0]+tmp[688]*kernel[1]+tmp[689]*kernel[2]+tmp[787]*kernel[3]+tmp[788]*kernel[4]+tmp[789]*kernel[5]+tmp[887]*kernel[6]+tmp[888]*kernel[7]+tmp[889]*kernel[8];
				ans[789]<=tmp[688]*kernel[0]+tmp[689]*kernel[1]+tmp[690]*kernel[2]+tmp[788]*kernel[3]+tmp[789]*kernel[4]+tmp[790]*kernel[5]+tmp[888]*kernel[6]+tmp[889]*kernel[7]+tmp[890]*kernel[8];
				ans[790]<=tmp[689]*kernel[0]+tmp[690]*kernel[1]+tmp[691]*kernel[2]+tmp[789]*kernel[3]+tmp[790]*kernel[4]+tmp[791]*kernel[5]+tmp[889]*kernel[6]+tmp[890]*kernel[7]+tmp[891]*kernel[8];
				ans[791]<=tmp[690]*kernel[0]+tmp[691]*kernel[1]+tmp[692]*kernel[2]+tmp[790]*kernel[3]+tmp[791]*kernel[4]+tmp[792]*kernel[5]+tmp[890]*kernel[6]+tmp[891]*kernel[7]+tmp[892]*kernel[8];
				ans[792]<=tmp[691]*kernel[0]+tmp[692]*kernel[1]+tmp[693]*kernel[2]+tmp[791]*kernel[3]+tmp[792]*kernel[4]+tmp[793]*kernel[5]+tmp[891]*kernel[6]+tmp[892]*kernel[7]+tmp[893]*kernel[8];
				ans[793]<=tmp[692]*kernel[0]+tmp[693]*kernel[1]+tmp[694]*kernel[2]+tmp[792]*kernel[3]+tmp[793]*kernel[4]+tmp[794]*kernel[5]+tmp[892]*kernel[6]+tmp[893]*kernel[7]+tmp[894]*kernel[8];
				ans[794]<=tmp[693]*kernel[0]+tmp[694]*kernel[1]+tmp[695]*kernel[2]+tmp[793]*kernel[3]+tmp[794]*kernel[4]+tmp[795]*kernel[5]+tmp[893]*kernel[6]+tmp[894]*kernel[7]+tmp[895]*kernel[8];
				ans[795]<=tmp[694]*kernel[0]+tmp[695]*kernel[1]+tmp[696]*kernel[2]+tmp[794]*kernel[3]+tmp[795]*kernel[4]+tmp[796]*kernel[5]+tmp[894]*kernel[6]+tmp[895]*kernel[7]+tmp[896]*kernel[8];
				ans[796]<=tmp[695]*kernel[0]+tmp[696]*kernel[1]+tmp[697]*kernel[2]+tmp[795]*kernel[3]+tmp[796]*kernel[4]+tmp[797]*kernel[5]+tmp[895]*kernel[6]+tmp[896]*kernel[7]+tmp[897]*kernel[8];
				ans[797]<=tmp[696]*kernel[0]+tmp[697]*kernel[1]+tmp[698]*kernel[2]+tmp[796]*kernel[3]+tmp[797]*kernel[4]+tmp[798]*kernel[5]+tmp[896]*kernel[6]+tmp[897]*kernel[7]+tmp[898]*kernel[8];
				ans[798]<=tmp[697]*kernel[0]+tmp[698]*kernel[1]+tmp[699]*kernel[2]+tmp[797]*kernel[3]+tmp[798]*kernel[4]+tmp[799]*kernel[5]+tmp[897]*kernel[6]+tmp[898]*kernel[7]+tmp[899]*kernel[8];
				ans[799]<=tmp[698]*kernel[0]+tmp[699]*kernel[1]+tmp[798]*kernel[3]+tmp[799]*kernel[4]+tmp[898]*kernel[6]+tmp[899]*kernel[7];
				ans[800]<=tmp[700]*kernel[1]+tmp[701]*kernel[2]+tmp[800]*kernel[4]+tmp[801]*kernel[5]+tmp[900]*kernel[7]+tmp[901]*kernel[8];
				ans[801]<=tmp[700]*kernel[0]+tmp[701]*kernel[1]+tmp[702]*kernel[2]+tmp[800]*kernel[3]+tmp[801]*kernel[4]+tmp[802]*kernel[5]+tmp[900]*kernel[6]+tmp[901]*kernel[7]+tmp[902]*kernel[8];
				ans[802]<=tmp[701]*kernel[0]+tmp[702]*kernel[1]+tmp[703]*kernel[2]+tmp[801]*kernel[3]+tmp[802]*kernel[4]+tmp[803]*kernel[5]+tmp[901]*kernel[6]+tmp[902]*kernel[7]+tmp[903]*kernel[8];
				ans[803]<=tmp[702]*kernel[0]+tmp[703]*kernel[1]+tmp[704]*kernel[2]+tmp[802]*kernel[3]+tmp[803]*kernel[4]+tmp[804]*kernel[5]+tmp[902]*kernel[6]+tmp[903]*kernel[7]+tmp[904]*kernel[8];
				ans[804]<=tmp[703]*kernel[0]+tmp[704]*kernel[1]+tmp[705]*kernel[2]+tmp[803]*kernel[3]+tmp[804]*kernel[4]+tmp[805]*kernel[5]+tmp[903]*kernel[6]+tmp[904]*kernel[7]+tmp[905]*kernel[8];
				ans[805]<=tmp[704]*kernel[0]+tmp[705]*kernel[1]+tmp[706]*kernel[2]+tmp[804]*kernel[3]+tmp[805]*kernel[4]+tmp[806]*kernel[5]+tmp[904]*kernel[6]+tmp[905]*kernel[7]+tmp[906]*kernel[8];
				ans[806]<=tmp[705]*kernel[0]+tmp[706]*kernel[1]+tmp[707]*kernel[2]+tmp[805]*kernel[3]+tmp[806]*kernel[4]+tmp[807]*kernel[5]+tmp[905]*kernel[6]+tmp[906]*kernel[7]+tmp[907]*kernel[8];
				ans[807]<=tmp[706]*kernel[0]+tmp[707]*kernel[1]+tmp[708]*kernel[2]+tmp[806]*kernel[3]+tmp[807]*kernel[4]+tmp[808]*kernel[5]+tmp[906]*kernel[6]+tmp[907]*kernel[7]+tmp[908]*kernel[8];
				ans[808]<=tmp[707]*kernel[0]+tmp[708]*kernel[1]+tmp[709]*kernel[2]+tmp[807]*kernel[3]+tmp[808]*kernel[4]+tmp[809]*kernel[5]+tmp[907]*kernel[6]+tmp[908]*kernel[7]+tmp[909]*kernel[8];
				ans[809]<=tmp[708]*kernel[0]+tmp[709]*kernel[1]+tmp[710]*kernel[2]+tmp[808]*kernel[3]+tmp[809]*kernel[4]+tmp[810]*kernel[5]+tmp[908]*kernel[6]+tmp[909]*kernel[7]+tmp[910]*kernel[8];
				ans[810]<=tmp[709]*kernel[0]+tmp[710]*kernel[1]+tmp[711]*kernel[2]+tmp[809]*kernel[3]+tmp[810]*kernel[4]+tmp[811]*kernel[5]+tmp[909]*kernel[6]+tmp[910]*kernel[7]+tmp[911]*kernel[8];
				ans[811]<=tmp[710]*kernel[0]+tmp[711]*kernel[1]+tmp[712]*kernel[2]+tmp[810]*kernel[3]+tmp[811]*kernel[4]+tmp[812]*kernel[5]+tmp[910]*kernel[6]+tmp[911]*kernel[7]+tmp[912]*kernel[8];
				ans[812]<=tmp[711]*kernel[0]+tmp[712]*kernel[1]+tmp[713]*kernel[2]+tmp[811]*kernel[3]+tmp[812]*kernel[4]+tmp[813]*kernel[5]+tmp[911]*kernel[6]+tmp[912]*kernel[7]+tmp[913]*kernel[8];
				ans[813]<=tmp[712]*kernel[0]+tmp[713]*kernel[1]+tmp[714]*kernel[2]+tmp[812]*kernel[3]+tmp[813]*kernel[4]+tmp[814]*kernel[5]+tmp[912]*kernel[6]+tmp[913]*kernel[7]+tmp[914]*kernel[8];
				ans[814]<=tmp[713]*kernel[0]+tmp[714]*kernel[1]+tmp[715]*kernel[2]+tmp[813]*kernel[3]+tmp[814]*kernel[4]+tmp[815]*kernel[5]+tmp[913]*kernel[6]+tmp[914]*kernel[7]+tmp[915]*kernel[8];
				ans[815]<=tmp[714]*kernel[0]+tmp[715]*kernel[1]+tmp[716]*kernel[2]+tmp[814]*kernel[3]+tmp[815]*kernel[4]+tmp[816]*kernel[5]+tmp[914]*kernel[6]+tmp[915]*kernel[7]+tmp[916]*kernel[8];
				ans[816]<=tmp[715]*kernel[0]+tmp[716]*kernel[1]+tmp[717]*kernel[2]+tmp[815]*kernel[3]+tmp[816]*kernel[4]+tmp[817]*kernel[5]+tmp[915]*kernel[6]+tmp[916]*kernel[7]+tmp[917]*kernel[8];
				ans[817]<=tmp[716]*kernel[0]+tmp[717]*kernel[1]+tmp[718]*kernel[2]+tmp[816]*kernel[3]+tmp[817]*kernel[4]+tmp[818]*kernel[5]+tmp[916]*kernel[6]+tmp[917]*kernel[7]+tmp[918]*kernel[8];
				ans[818]<=tmp[717]*kernel[0]+tmp[718]*kernel[1]+tmp[719]*kernel[2]+tmp[817]*kernel[3]+tmp[818]*kernel[4]+tmp[819]*kernel[5]+tmp[917]*kernel[6]+tmp[918]*kernel[7]+tmp[919]*kernel[8];
				ans[819]<=tmp[718]*kernel[0]+tmp[719]*kernel[1]+tmp[720]*kernel[2]+tmp[818]*kernel[3]+tmp[819]*kernel[4]+tmp[820]*kernel[5]+tmp[918]*kernel[6]+tmp[919]*kernel[7]+tmp[920]*kernel[8];
				ans[820]<=tmp[719]*kernel[0]+tmp[720]*kernel[1]+tmp[721]*kernel[2]+tmp[819]*kernel[3]+tmp[820]*kernel[4]+tmp[821]*kernel[5]+tmp[919]*kernel[6]+tmp[920]*kernel[7]+tmp[921]*kernel[8];
				ans[821]<=tmp[720]*kernel[0]+tmp[721]*kernel[1]+tmp[722]*kernel[2]+tmp[820]*kernel[3]+tmp[821]*kernel[4]+tmp[822]*kernel[5]+tmp[920]*kernel[6]+tmp[921]*kernel[7]+tmp[922]*kernel[8];
				ans[822]<=tmp[721]*kernel[0]+tmp[722]*kernel[1]+tmp[723]*kernel[2]+tmp[821]*kernel[3]+tmp[822]*kernel[4]+tmp[823]*kernel[5]+tmp[921]*kernel[6]+tmp[922]*kernel[7]+tmp[923]*kernel[8];
				ans[823]<=tmp[722]*kernel[0]+tmp[723]*kernel[1]+tmp[724]*kernel[2]+tmp[822]*kernel[3]+tmp[823]*kernel[4]+tmp[824]*kernel[5]+tmp[922]*kernel[6]+tmp[923]*kernel[7]+tmp[924]*kernel[8];
				ans[824]<=tmp[723]*kernel[0]+tmp[724]*kernel[1]+tmp[725]*kernel[2]+tmp[823]*kernel[3]+tmp[824]*kernel[4]+tmp[825]*kernel[5]+tmp[923]*kernel[6]+tmp[924]*kernel[7]+tmp[925]*kernel[8];
				ans[825]<=tmp[724]*kernel[0]+tmp[725]*kernel[1]+tmp[726]*kernel[2]+tmp[824]*kernel[3]+tmp[825]*kernel[4]+tmp[826]*kernel[5]+tmp[924]*kernel[6]+tmp[925]*kernel[7]+tmp[926]*kernel[8];
				ans[826]<=tmp[725]*kernel[0]+tmp[726]*kernel[1]+tmp[727]*kernel[2]+tmp[825]*kernel[3]+tmp[826]*kernel[4]+tmp[827]*kernel[5]+tmp[925]*kernel[6]+tmp[926]*kernel[7]+tmp[927]*kernel[8];
				ans[827]<=tmp[726]*kernel[0]+tmp[727]*kernel[1]+tmp[728]*kernel[2]+tmp[826]*kernel[3]+tmp[827]*kernel[4]+tmp[828]*kernel[5]+tmp[926]*kernel[6]+tmp[927]*kernel[7]+tmp[928]*kernel[8];
				ans[828]<=tmp[727]*kernel[0]+tmp[728]*kernel[1]+tmp[729]*kernel[2]+tmp[827]*kernel[3]+tmp[828]*kernel[4]+tmp[829]*kernel[5]+tmp[927]*kernel[6]+tmp[928]*kernel[7]+tmp[929]*kernel[8];
				ans[829]<=tmp[728]*kernel[0]+tmp[729]*kernel[1]+tmp[730]*kernel[2]+tmp[828]*kernel[3]+tmp[829]*kernel[4]+tmp[830]*kernel[5]+tmp[928]*kernel[6]+tmp[929]*kernel[7]+tmp[930]*kernel[8];
				ans[830]<=tmp[729]*kernel[0]+tmp[730]*kernel[1]+tmp[731]*kernel[2]+tmp[829]*kernel[3]+tmp[830]*kernel[4]+tmp[831]*kernel[5]+tmp[929]*kernel[6]+tmp[930]*kernel[7]+tmp[931]*kernel[8];
				ans[831]<=tmp[730]*kernel[0]+tmp[731]*kernel[1]+tmp[732]*kernel[2]+tmp[830]*kernel[3]+tmp[831]*kernel[4]+tmp[832]*kernel[5]+tmp[930]*kernel[6]+tmp[931]*kernel[7]+tmp[932]*kernel[8];
				ans[832]<=tmp[731]*kernel[0]+tmp[732]*kernel[1]+tmp[733]*kernel[2]+tmp[831]*kernel[3]+tmp[832]*kernel[4]+tmp[833]*kernel[5]+tmp[931]*kernel[6]+tmp[932]*kernel[7]+tmp[933]*kernel[8];
				ans[833]<=tmp[732]*kernel[0]+tmp[733]*kernel[1]+tmp[734]*kernel[2]+tmp[832]*kernel[3]+tmp[833]*kernel[4]+tmp[834]*kernel[5]+tmp[932]*kernel[6]+tmp[933]*kernel[7]+tmp[934]*kernel[8];
				ans[834]<=tmp[733]*kernel[0]+tmp[734]*kernel[1]+tmp[735]*kernel[2]+tmp[833]*kernel[3]+tmp[834]*kernel[4]+tmp[835]*kernel[5]+tmp[933]*kernel[6]+tmp[934]*kernel[7]+tmp[935]*kernel[8];
				ans[835]<=tmp[734]*kernel[0]+tmp[735]*kernel[1]+tmp[736]*kernel[2]+tmp[834]*kernel[3]+tmp[835]*kernel[4]+tmp[836]*kernel[5]+tmp[934]*kernel[6]+tmp[935]*kernel[7]+tmp[936]*kernel[8];
				ans[836]<=tmp[735]*kernel[0]+tmp[736]*kernel[1]+tmp[737]*kernel[2]+tmp[835]*kernel[3]+tmp[836]*kernel[4]+tmp[837]*kernel[5]+tmp[935]*kernel[6]+tmp[936]*kernel[7]+tmp[937]*kernel[8];
				ans[837]<=tmp[736]*kernel[0]+tmp[737]*kernel[1]+tmp[738]*kernel[2]+tmp[836]*kernel[3]+tmp[837]*kernel[4]+tmp[838]*kernel[5]+tmp[936]*kernel[6]+tmp[937]*kernel[7]+tmp[938]*kernel[8];
				ans[838]<=tmp[737]*kernel[0]+tmp[738]*kernel[1]+tmp[739]*kernel[2]+tmp[837]*kernel[3]+tmp[838]*kernel[4]+tmp[839]*kernel[5]+tmp[937]*kernel[6]+tmp[938]*kernel[7]+tmp[939]*kernel[8];
				ans[839]<=tmp[738]*kernel[0]+tmp[739]*kernel[1]+tmp[740]*kernel[2]+tmp[838]*kernel[3]+tmp[839]*kernel[4]+tmp[840]*kernel[5]+tmp[938]*kernel[6]+tmp[939]*kernel[7]+tmp[940]*kernel[8];
				ans[840]<=tmp[739]*kernel[0]+tmp[740]*kernel[1]+tmp[741]*kernel[2]+tmp[839]*kernel[3]+tmp[840]*kernel[4]+tmp[841]*kernel[5]+tmp[939]*kernel[6]+tmp[940]*kernel[7]+tmp[941]*kernel[8];
				ans[841]<=tmp[740]*kernel[0]+tmp[741]*kernel[1]+tmp[742]*kernel[2]+tmp[840]*kernel[3]+tmp[841]*kernel[4]+tmp[842]*kernel[5]+tmp[940]*kernel[6]+tmp[941]*kernel[7]+tmp[942]*kernel[8];
				ans[842]<=tmp[741]*kernel[0]+tmp[742]*kernel[1]+tmp[743]*kernel[2]+tmp[841]*kernel[3]+tmp[842]*kernel[4]+tmp[843]*kernel[5]+tmp[941]*kernel[6]+tmp[942]*kernel[7]+tmp[943]*kernel[8];
				ans[843]<=tmp[742]*kernel[0]+tmp[743]*kernel[1]+tmp[744]*kernel[2]+tmp[842]*kernel[3]+tmp[843]*kernel[4]+tmp[844]*kernel[5]+tmp[942]*kernel[6]+tmp[943]*kernel[7]+tmp[944]*kernel[8];
				ans[844]<=tmp[743]*kernel[0]+tmp[744]*kernel[1]+tmp[745]*kernel[2]+tmp[843]*kernel[3]+tmp[844]*kernel[4]+tmp[845]*kernel[5]+tmp[943]*kernel[6]+tmp[944]*kernel[7]+tmp[945]*kernel[8];
				ans[845]<=tmp[744]*kernel[0]+tmp[745]*kernel[1]+tmp[746]*kernel[2]+tmp[844]*kernel[3]+tmp[845]*kernel[4]+tmp[846]*kernel[5]+tmp[944]*kernel[6]+tmp[945]*kernel[7]+tmp[946]*kernel[8];
				ans[846]<=tmp[745]*kernel[0]+tmp[746]*kernel[1]+tmp[747]*kernel[2]+tmp[845]*kernel[3]+tmp[846]*kernel[4]+tmp[847]*kernel[5]+tmp[945]*kernel[6]+tmp[946]*kernel[7]+tmp[947]*kernel[8];
				ans[847]<=tmp[746]*kernel[0]+tmp[747]*kernel[1]+tmp[748]*kernel[2]+tmp[846]*kernel[3]+tmp[847]*kernel[4]+tmp[848]*kernel[5]+tmp[946]*kernel[6]+tmp[947]*kernel[7]+tmp[948]*kernel[8];
				ans[848]<=tmp[747]*kernel[0]+tmp[748]*kernel[1]+tmp[749]*kernel[2]+tmp[847]*kernel[3]+tmp[848]*kernel[4]+tmp[849]*kernel[5]+tmp[947]*kernel[6]+tmp[948]*kernel[7]+tmp[949]*kernel[8];
				ans[849]<=tmp[748]*kernel[0]+tmp[749]*kernel[1]+tmp[750]*kernel[2]+tmp[848]*kernel[3]+tmp[849]*kernel[4]+tmp[850]*kernel[5]+tmp[948]*kernel[6]+tmp[949]*kernel[7]+tmp[950]*kernel[8];
				ans[850]<=tmp[749]*kernel[0]+tmp[750]*kernel[1]+tmp[751]*kernel[2]+tmp[849]*kernel[3]+tmp[850]*kernel[4]+tmp[851]*kernel[5]+tmp[949]*kernel[6]+tmp[950]*kernel[7]+tmp[951]*kernel[8];
				ans[851]<=tmp[750]*kernel[0]+tmp[751]*kernel[1]+tmp[752]*kernel[2]+tmp[850]*kernel[3]+tmp[851]*kernel[4]+tmp[852]*kernel[5]+tmp[950]*kernel[6]+tmp[951]*kernel[7]+tmp[952]*kernel[8];
				ans[852]<=tmp[751]*kernel[0]+tmp[752]*kernel[1]+tmp[753]*kernel[2]+tmp[851]*kernel[3]+tmp[852]*kernel[4]+tmp[853]*kernel[5]+tmp[951]*kernel[6]+tmp[952]*kernel[7]+tmp[953]*kernel[8];
				ans[853]<=tmp[752]*kernel[0]+tmp[753]*kernel[1]+tmp[754]*kernel[2]+tmp[852]*kernel[3]+tmp[853]*kernel[4]+tmp[854]*kernel[5]+tmp[952]*kernel[6]+tmp[953]*kernel[7]+tmp[954]*kernel[8];
				ans[854]<=tmp[753]*kernel[0]+tmp[754]*kernel[1]+tmp[755]*kernel[2]+tmp[853]*kernel[3]+tmp[854]*kernel[4]+tmp[855]*kernel[5]+tmp[953]*kernel[6]+tmp[954]*kernel[7]+tmp[955]*kernel[8];
				ans[855]<=tmp[754]*kernel[0]+tmp[755]*kernel[1]+tmp[756]*kernel[2]+tmp[854]*kernel[3]+tmp[855]*kernel[4]+tmp[856]*kernel[5]+tmp[954]*kernel[6]+tmp[955]*kernel[7]+tmp[956]*kernel[8];
				ans[856]<=tmp[755]*kernel[0]+tmp[756]*kernel[1]+tmp[757]*kernel[2]+tmp[855]*kernel[3]+tmp[856]*kernel[4]+tmp[857]*kernel[5]+tmp[955]*kernel[6]+tmp[956]*kernel[7]+tmp[957]*kernel[8];
				ans[857]<=tmp[756]*kernel[0]+tmp[757]*kernel[1]+tmp[758]*kernel[2]+tmp[856]*kernel[3]+tmp[857]*kernel[4]+tmp[858]*kernel[5]+tmp[956]*kernel[6]+tmp[957]*kernel[7]+tmp[958]*kernel[8];
				ans[858]<=tmp[757]*kernel[0]+tmp[758]*kernel[1]+tmp[759]*kernel[2]+tmp[857]*kernel[3]+tmp[858]*kernel[4]+tmp[859]*kernel[5]+tmp[957]*kernel[6]+tmp[958]*kernel[7]+tmp[959]*kernel[8];
				ans[859]<=tmp[758]*kernel[0]+tmp[759]*kernel[1]+tmp[760]*kernel[2]+tmp[858]*kernel[3]+tmp[859]*kernel[4]+tmp[860]*kernel[5]+tmp[958]*kernel[6]+tmp[959]*kernel[7]+tmp[960]*kernel[8];
				ans[860]<=tmp[759]*kernel[0]+tmp[760]*kernel[1]+tmp[761]*kernel[2]+tmp[859]*kernel[3]+tmp[860]*kernel[4]+tmp[861]*kernel[5]+tmp[959]*kernel[6]+tmp[960]*kernel[7]+tmp[961]*kernel[8];
				ans[861]<=tmp[760]*kernel[0]+tmp[761]*kernel[1]+tmp[762]*kernel[2]+tmp[860]*kernel[3]+tmp[861]*kernel[4]+tmp[862]*kernel[5]+tmp[960]*kernel[6]+tmp[961]*kernel[7]+tmp[962]*kernel[8];
				ans[862]<=tmp[761]*kernel[0]+tmp[762]*kernel[1]+tmp[763]*kernel[2]+tmp[861]*kernel[3]+tmp[862]*kernel[4]+tmp[863]*kernel[5]+tmp[961]*kernel[6]+tmp[962]*kernel[7]+tmp[963]*kernel[8];
				ans[863]<=tmp[762]*kernel[0]+tmp[763]*kernel[1]+tmp[764]*kernel[2]+tmp[862]*kernel[3]+tmp[863]*kernel[4]+tmp[864]*kernel[5]+tmp[962]*kernel[6]+tmp[963]*kernel[7]+tmp[964]*kernel[8];
				ans[864]<=tmp[763]*kernel[0]+tmp[764]*kernel[1]+tmp[765]*kernel[2]+tmp[863]*kernel[3]+tmp[864]*kernel[4]+tmp[865]*kernel[5]+tmp[963]*kernel[6]+tmp[964]*kernel[7]+tmp[965]*kernel[8];
				ans[865]<=tmp[764]*kernel[0]+tmp[765]*kernel[1]+tmp[766]*kernel[2]+tmp[864]*kernel[3]+tmp[865]*kernel[4]+tmp[866]*kernel[5]+tmp[964]*kernel[6]+tmp[965]*kernel[7]+tmp[966]*kernel[8];
				ans[866]<=tmp[765]*kernel[0]+tmp[766]*kernel[1]+tmp[767]*kernel[2]+tmp[865]*kernel[3]+tmp[866]*kernel[4]+tmp[867]*kernel[5]+tmp[965]*kernel[6]+tmp[966]*kernel[7]+tmp[967]*kernel[8];
				ans[867]<=tmp[766]*kernel[0]+tmp[767]*kernel[1]+tmp[768]*kernel[2]+tmp[866]*kernel[3]+tmp[867]*kernel[4]+tmp[868]*kernel[5]+tmp[966]*kernel[6]+tmp[967]*kernel[7]+tmp[968]*kernel[8];
				ans[868]<=tmp[767]*kernel[0]+tmp[768]*kernel[1]+tmp[769]*kernel[2]+tmp[867]*kernel[3]+tmp[868]*kernel[4]+tmp[869]*kernel[5]+tmp[967]*kernel[6]+tmp[968]*kernel[7]+tmp[969]*kernel[8];
				ans[869]<=tmp[768]*kernel[0]+tmp[769]*kernel[1]+tmp[770]*kernel[2]+tmp[868]*kernel[3]+tmp[869]*kernel[4]+tmp[870]*kernel[5]+tmp[968]*kernel[6]+tmp[969]*kernel[7]+tmp[970]*kernel[8];
				ans[870]<=tmp[769]*kernel[0]+tmp[770]*kernel[1]+tmp[771]*kernel[2]+tmp[869]*kernel[3]+tmp[870]*kernel[4]+tmp[871]*kernel[5]+tmp[969]*kernel[6]+tmp[970]*kernel[7]+tmp[971]*kernel[8];
				ans[871]<=tmp[770]*kernel[0]+tmp[771]*kernel[1]+tmp[772]*kernel[2]+tmp[870]*kernel[3]+tmp[871]*kernel[4]+tmp[872]*kernel[5]+tmp[970]*kernel[6]+tmp[971]*kernel[7]+tmp[972]*kernel[8];
				ans[872]<=tmp[771]*kernel[0]+tmp[772]*kernel[1]+tmp[773]*kernel[2]+tmp[871]*kernel[3]+tmp[872]*kernel[4]+tmp[873]*kernel[5]+tmp[971]*kernel[6]+tmp[972]*kernel[7]+tmp[973]*kernel[8];
				ans[873]<=tmp[772]*kernel[0]+tmp[773]*kernel[1]+tmp[774]*kernel[2]+tmp[872]*kernel[3]+tmp[873]*kernel[4]+tmp[874]*kernel[5]+tmp[972]*kernel[6]+tmp[973]*kernel[7]+tmp[974]*kernel[8];
				ans[874]<=tmp[773]*kernel[0]+tmp[774]*kernel[1]+tmp[775]*kernel[2]+tmp[873]*kernel[3]+tmp[874]*kernel[4]+tmp[875]*kernel[5]+tmp[973]*kernel[6]+tmp[974]*kernel[7]+tmp[975]*kernel[8];
				ans[875]<=tmp[774]*kernel[0]+tmp[775]*kernel[1]+tmp[776]*kernel[2]+tmp[874]*kernel[3]+tmp[875]*kernel[4]+tmp[876]*kernel[5]+tmp[974]*kernel[6]+tmp[975]*kernel[7]+tmp[976]*kernel[8];
				ans[876]<=tmp[775]*kernel[0]+tmp[776]*kernel[1]+tmp[777]*kernel[2]+tmp[875]*kernel[3]+tmp[876]*kernel[4]+tmp[877]*kernel[5]+tmp[975]*kernel[6]+tmp[976]*kernel[7]+tmp[977]*kernel[8];
				ans[877]<=tmp[776]*kernel[0]+tmp[777]*kernel[1]+tmp[778]*kernel[2]+tmp[876]*kernel[3]+tmp[877]*kernel[4]+tmp[878]*kernel[5]+tmp[976]*kernel[6]+tmp[977]*kernel[7]+tmp[978]*kernel[8];
				ans[878]<=tmp[777]*kernel[0]+tmp[778]*kernel[1]+tmp[779]*kernel[2]+tmp[877]*kernel[3]+tmp[878]*kernel[4]+tmp[879]*kernel[5]+tmp[977]*kernel[6]+tmp[978]*kernel[7]+tmp[979]*kernel[8];
				ans[879]<=tmp[778]*kernel[0]+tmp[779]*kernel[1]+tmp[780]*kernel[2]+tmp[878]*kernel[3]+tmp[879]*kernel[4]+tmp[880]*kernel[5]+tmp[978]*kernel[6]+tmp[979]*kernel[7]+tmp[980]*kernel[8];
				ans[880]<=tmp[779]*kernel[0]+tmp[780]*kernel[1]+tmp[781]*kernel[2]+tmp[879]*kernel[3]+tmp[880]*kernel[4]+tmp[881]*kernel[5]+tmp[979]*kernel[6]+tmp[980]*kernel[7]+tmp[981]*kernel[8];
				ans[881]<=tmp[780]*kernel[0]+tmp[781]*kernel[1]+tmp[782]*kernel[2]+tmp[880]*kernel[3]+tmp[881]*kernel[4]+tmp[882]*kernel[5]+tmp[980]*kernel[6]+tmp[981]*kernel[7]+tmp[982]*kernel[8];
				ans[882]<=tmp[781]*kernel[0]+tmp[782]*kernel[1]+tmp[783]*kernel[2]+tmp[881]*kernel[3]+tmp[882]*kernel[4]+tmp[883]*kernel[5]+tmp[981]*kernel[6]+tmp[982]*kernel[7]+tmp[983]*kernel[8];
				ans[883]<=tmp[782]*kernel[0]+tmp[783]*kernel[1]+tmp[784]*kernel[2]+tmp[882]*kernel[3]+tmp[883]*kernel[4]+tmp[884]*kernel[5]+tmp[982]*kernel[6]+tmp[983]*kernel[7]+tmp[984]*kernel[8];
				ans[884]<=tmp[783]*kernel[0]+tmp[784]*kernel[1]+tmp[785]*kernel[2]+tmp[883]*kernel[3]+tmp[884]*kernel[4]+tmp[885]*kernel[5]+tmp[983]*kernel[6]+tmp[984]*kernel[7]+tmp[985]*kernel[8];
				ans[885]<=tmp[784]*kernel[0]+tmp[785]*kernel[1]+tmp[786]*kernel[2]+tmp[884]*kernel[3]+tmp[885]*kernel[4]+tmp[886]*kernel[5]+tmp[984]*kernel[6]+tmp[985]*kernel[7]+tmp[986]*kernel[8];
				ans[886]<=tmp[785]*kernel[0]+tmp[786]*kernel[1]+tmp[787]*kernel[2]+tmp[885]*kernel[3]+tmp[886]*kernel[4]+tmp[887]*kernel[5]+tmp[985]*kernel[6]+tmp[986]*kernel[7]+tmp[987]*kernel[8];
				ans[887]<=tmp[786]*kernel[0]+tmp[787]*kernel[1]+tmp[788]*kernel[2]+tmp[886]*kernel[3]+tmp[887]*kernel[4]+tmp[888]*kernel[5]+tmp[986]*kernel[6]+tmp[987]*kernel[7]+tmp[988]*kernel[8];
				ans[888]<=tmp[787]*kernel[0]+tmp[788]*kernel[1]+tmp[789]*kernel[2]+tmp[887]*kernel[3]+tmp[888]*kernel[4]+tmp[889]*kernel[5]+tmp[987]*kernel[6]+tmp[988]*kernel[7]+tmp[989]*kernel[8];
				ans[889]<=tmp[788]*kernel[0]+tmp[789]*kernel[1]+tmp[790]*kernel[2]+tmp[888]*kernel[3]+tmp[889]*kernel[4]+tmp[890]*kernel[5]+tmp[988]*kernel[6]+tmp[989]*kernel[7]+tmp[990]*kernel[8];
				ans[890]<=tmp[789]*kernel[0]+tmp[790]*kernel[1]+tmp[791]*kernel[2]+tmp[889]*kernel[3]+tmp[890]*kernel[4]+tmp[891]*kernel[5]+tmp[989]*kernel[6]+tmp[990]*kernel[7]+tmp[991]*kernel[8];
				ans[891]<=tmp[790]*kernel[0]+tmp[791]*kernel[1]+tmp[792]*kernel[2]+tmp[890]*kernel[3]+tmp[891]*kernel[4]+tmp[892]*kernel[5]+tmp[990]*kernel[6]+tmp[991]*kernel[7]+tmp[992]*kernel[8];
				ans[892]<=tmp[791]*kernel[0]+tmp[792]*kernel[1]+tmp[793]*kernel[2]+tmp[891]*kernel[3]+tmp[892]*kernel[4]+tmp[893]*kernel[5]+tmp[991]*kernel[6]+tmp[992]*kernel[7]+tmp[993]*kernel[8];
				ans[893]<=tmp[792]*kernel[0]+tmp[793]*kernel[1]+tmp[794]*kernel[2]+tmp[892]*kernel[3]+tmp[893]*kernel[4]+tmp[894]*kernel[5]+tmp[992]*kernel[6]+tmp[993]*kernel[7]+tmp[994]*kernel[8];
				ans[894]<=tmp[793]*kernel[0]+tmp[794]*kernel[1]+tmp[795]*kernel[2]+tmp[893]*kernel[3]+tmp[894]*kernel[4]+tmp[895]*kernel[5]+tmp[993]*kernel[6]+tmp[994]*kernel[7]+tmp[995]*kernel[8];
				ans[895]<=tmp[794]*kernel[0]+tmp[795]*kernel[1]+tmp[796]*kernel[2]+tmp[894]*kernel[3]+tmp[895]*kernel[4]+tmp[896]*kernel[5]+tmp[994]*kernel[6]+tmp[995]*kernel[7]+tmp[996]*kernel[8];
				ans[896]<=tmp[795]*kernel[0]+tmp[796]*kernel[1]+tmp[797]*kernel[2]+tmp[895]*kernel[3]+tmp[896]*kernel[4]+tmp[897]*kernel[5]+tmp[995]*kernel[6]+tmp[996]*kernel[7]+tmp[997]*kernel[8];
				ans[897]<=tmp[796]*kernel[0]+tmp[797]*kernel[1]+tmp[798]*kernel[2]+tmp[896]*kernel[3]+tmp[897]*kernel[4]+tmp[898]*kernel[5]+tmp[996]*kernel[6]+tmp[997]*kernel[7]+tmp[998]*kernel[8];
				ans[898]<=tmp[797]*kernel[0]+tmp[798]*kernel[1]+tmp[799]*kernel[2]+tmp[897]*kernel[3]+tmp[898]*kernel[4]+tmp[899]*kernel[5]+tmp[997]*kernel[6]+tmp[998]*kernel[7]+tmp[999]*kernel[8];
				ans[899]<=tmp[798]*kernel[0]+tmp[799]*kernel[1]+tmp[898]*kernel[3]+tmp[899]*kernel[4]+tmp[998]*kernel[6]+tmp[999]*kernel[7];
				ans[900]<=tmp[800]*kernel[1]+tmp[801]*kernel[2]+tmp[900]*kernel[4]+tmp[901]*kernel[5]+tmp[1000]*kernel[7]+tmp[1001]*kernel[8];
				ans[901]<=tmp[800]*kernel[0]+tmp[801]*kernel[1]+tmp[802]*kernel[2]+tmp[900]*kernel[3]+tmp[901]*kernel[4]+tmp[902]*kernel[5]+tmp[1000]*kernel[6]+tmp[1001]*kernel[7]+tmp[1002]*kernel[8];
				ans[902]<=tmp[801]*kernel[0]+tmp[802]*kernel[1]+tmp[803]*kernel[2]+tmp[901]*kernel[3]+tmp[902]*kernel[4]+tmp[903]*kernel[5]+tmp[1001]*kernel[6]+tmp[1002]*kernel[7]+tmp[1003]*kernel[8];
				ans[903]<=tmp[802]*kernel[0]+tmp[803]*kernel[1]+tmp[804]*kernel[2]+tmp[902]*kernel[3]+tmp[903]*kernel[4]+tmp[904]*kernel[5]+tmp[1002]*kernel[6]+tmp[1003]*kernel[7]+tmp[1004]*kernel[8];
				ans[904]<=tmp[803]*kernel[0]+tmp[804]*kernel[1]+tmp[805]*kernel[2]+tmp[903]*kernel[3]+tmp[904]*kernel[4]+tmp[905]*kernel[5]+tmp[1003]*kernel[6]+tmp[1004]*kernel[7]+tmp[1005]*kernel[8];
				ans[905]<=tmp[804]*kernel[0]+tmp[805]*kernel[1]+tmp[806]*kernel[2]+tmp[904]*kernel[3]+tmp[905]*kernel[4]+tmp[906]*kernel[5]+tmp[1004]*kernel[6]+tmp[1005]*kernel[7]+tmp[1006]*kernel[8];
				ans[906]<=tmp[805]*kernel[0]+tmp[806]*kernel[1]+tmp[807]*kernel[2]+tmp[905]*kernel[3]+tmp[906]*kernel[4]+tmp[907]*kernel[5]+tmp[1005]*kernel[6]+tmp[1006]*kernel[7]+tmp[1007]*kernel[8];
				ans[907]<=tmp[806]*kernel[0]+tmp[807]*kernel[1]+tmp[808]*kernel[2]+tmp[906]*kernel[3]+tmp[907]*kernel[4]+tmp[908]*kernel[5]+tmp[1006]*kernel[6]+tmp[1007]*kernel[7]+tmp[1008]*kernel[8];
				ans[908]<=tmp[807]*kernel[0]+tmp[808]*kernel[1]+tmp[809]*kernel[2]+tmp[907]*kernel[3]+tmp[908]*kernel[4]+tmp[909]*kernel[5]+tmp[1007]*kernel[6]+tmp[1008]*kernel[7]+tmp[1009]*kernel[8];
				ans[909]<=tmp[808]*kernel[0]+tmp[809]*kernel[1]+tmp[810]*kernel[2]+tmp[908]*kernel[3]+tmp[909]*kernel[4]+tmp[910]*kernel[5]+tmp[1008]*kernel[6]+tmp[1009]*kernel[7]+tmp[1010]*kernel[8];
				ans[910]<=tmp[809]*kernel[0]+tmp[810]*kernel[1]+tmp[811]*kernel[2]+tmp[909]*kernel[3]+tmp[910]*kernel[4]+tmp[911]*kernel[5]+tmp[1009]*kernel[6]+tmp[1010]*kernel[7]+tmp[1011]*kernel[8];
				ans[911]<=tmp[810]*kernel[0]+tmp[811]*kernel[1]+tmp[812]*kernel[2]+tmp[910]*kernel[3]+tmp[911]*kernel[4]+tmp[912]*kernel[5]+tmp[1010]*kernel[6]+tmp[1011]*kernel[7]+tmp[1012]*kernel[8];
				ans[912]<=tmp[811]*kernel[0]+tmp[812]*kernel[1]+tmp[813]*kernel[2]+tmp[911]*kernel[3]+tmp[912]*kernel[4]+tmp[913]*kernel[5]+tmp[1011]*kernel[6]+tmp[1012]*kernel[7]+tmp[1013]*kernel[8];
				ans[913]<=tmp[812]*kernel[0]+tmp[813]*kernel[1]+tmp[814]*kernel[2]+tmp[912]*kernel[3]+tmp[913]*kernel[4]+tmp[914]*kernel[5]+tmp[1012]*kernel[6]+tmp[1013]*kernel[7]+tmp[1014]*kernel[8];
				ans[914]<=tmp[813]*kernel[0]+tmp[814]*kernel[1]+tmp[815]*kernel[2]+tmp[913]*kernel[3]+tmp[914]*kernel[4]+tmp[915]*kernel[5]+tmp[1013]*kernel[6]+tmp[1014]*kernel[7]+tmp[1015]*kernel[8];
				ans[915]<=tmp[814]*kernel[0]+tmp[815]*kernel[1]+tmp[816]*kernel[2]+tmp[914]*kernel[3]+tmp[915]*kernel[4]+tmp[916]*kernel[5]+tmp[1014]*kernel[6]+tmp[1015]*kernel[7]+tmp[1016]*kernel[8];
				ans[916]<=tmp[815]*kernel[0]+tmp[816]*kernel[1]+tmp[817]*kernel[2]+tmp[915]*kernel[3]+tmp[916]*kernel[4]+tmp[917]*kernel[5]+tmp[1015]*kernel[6]+tmp[1016]*kernel[7]+tmp[1017]*kernel[8];
				ans[917]<=tmp[816]*kernel[0]+tmp[817]*kernel[1]+tmp[818]*kernel[2]+tmp[916]*kernel[3]+tmp[917]*kernel[4]+tmp[918]*kernel[5]+tmp[1016]*kernel[6]+tmp[1017]*kernel[7]+tmp[1018]*kernel[8];
				ans[918]<=tmp[817]*kernel[0]+tmp[818]*kernel[1]+tmp[819]*kernel[2]+tmp[917]*kernel[3]+tmp[918]*kernel[4]+tmp[919]*kernel[5]+tmp[1017]*kernel[6]+tmp[1018]*kernel[7]+tmp[1019]*kernel[8];
				ans[919]<=tmp[818]*kernel[0]+tmp[819]*kernel[1]+tmp[820]*kernel[2]+tmp[918]*kernel[3]+tmp[919]*kernel[4]+tmp[920]*kernel[5]+tmp[1018]*kernel[6]+tmp[1019]*kernel[7]+tmp[1020]*kernel[8];
				ans[920]<=tmp[819]*kernel[0]+tmp[820]*kernel[1]+tmp[821]*kernel[2]+tmp[919]*kernel[3]+tmp[920]*kernel[4]+tmp[921]*kernel[5]+tmp[1019]*kernel[6]+tmp[1020]*kernel[7]+tmp[1021]*kernel[8];
				ans[921]<=tmp[820]*kernel[0]+tmp[821]*kernel[1]+tmp[822]*kernel[2]+tmp[920]*kernel[3]+tmp[921]*kernel[4]+tmp[922]*kernel[5]+tmp[1020]*kernel[6]+tmp[1021]*kernel[7]+tmp[1022]*kernel[8];
				ans[922]<=tmp[821]*kernel[0]+tmp[822]*kernel[1]+tmp[823]*kernel[2]+tmp[921]*kernel[3]+tmp[922]*kernel[4]+tmp[923]*kernel[5]+tmp[1021]*kernel[6]+tmp[1022]*kernel[7]+tmp[1023]*kernel[8];
				ans[923]<=tmp[822]*kernel[0]+tmp[823]*kernel[1]+tmp[824]*kernel[2]+tmp[922]*kernel[3]+tmp[923]*kernel[4]+tmp[924]*kernel[5]+tmp[1022]*kernel[6]+tmp[1023]*kernel[7]+tmp[1024]*kernel[8];
				ans[924]<=tmp[823]*kernel[0]+tmp[824]*kernel[1]+tmp[825]*kernel[2]+tmp[923]*kernel[3]+tmp[924]*kernel[4]+tmp[925]*kernel[5]+tmp[1023]*kernel[6]+tmp[1024]*kernel[7]+tmp[1025]*kernel[8];
				ans[925]<=tmp[824]*kernel[0]+tmp[825]*kernel[1]+tmp[826]*kernel[2]+tmp[924]*kernel[3]+tmp[925]*kernel[4]+tmp[926]*kernel[5]+tmp[1024]*kernel[6]+tmp[1025]*kernel[7]+tmp[1026]*kernel[8];
				ans[926]<=tmp[825]*kernel[0]+tmp[826]*kernel[1]+tmp[827]*kernel[2]+tmp[925]*kernel[3]+tmp[926]*kernel[4]+tmp[927]*kernel[5]+tmp[1025]*kernel[6]+tmp[1026]*kernel[7]+tmp[1027]*kernel[8];
				ans[927]<=tmp[826]*kernel[0]+tmp[827]*kernel[1]+tmp[828]*kernel[2]+tmp[926]*kernel[3]+tmp[927]*kernel[4]+tmp[928]*kernel[5]+tmp[1026]*kernel[6]+tmp[1027]*kernel[7]+tmp[1028]*kernel[8];
				ans[928]<=tmp[827]*kernel[0]+tmp[828]*kernel[1]+tmp[829]*kernel[2]+tmp[927]*kernel[3]+tmp[928]*kernel[4]+tmp[929]*kernel[5]+tmp[1027]*kernel[6]+tmp[1028]*kernel[7]+tmp[1029]*kernel[8];
				ans[929]<=tmp[828]*kernel[0]+tmp[829]*kernel[1]+tmp[830]*kernel[2]+tmp[928]*kernel[3]+tmp[929]*kernel[4]+tmp[930]*kernel[5]+tmp[1028]*kernel[6]+tmp[1029]*kernel[7]+tmp[1030]*kernel[8];
				ans[930]<=tmp[829]*kernel[0]+tmp[830]*kernel[1]+tmp[831]*kernel[2]+tmp[929]*kernel[3]+tmp[930]*kernel[4]+tmp[931]*kernel[5]+tmp[1029]*kernel[6]+tmp[1030]*kernel[7]+tmp[1031]*kernel[8];
				ans[931]<=tmp[830]*kernel[0]+tmp[831]*kernel[1]+tmp[832]*kernel[2]+tmp[930]*kernel[3]+tmp[931]*kernel[4]+tmp[932]*kernel[5]+tmp[1030]*kernel[6]+tmp[1031]*kernel[7]+tmp[1032]*kernel[8];
				ans[932]<=tmp[831]*kernel[0]+tmp[832]*kernel[1]+tmp[833]*kernel[2]+tmp[931]*kernel[3]+tmp[932]*kernel[4]+tmp[933]*kernel[5]+tmp[1031]*kernel[6]+tmp[1032]*kernel[7]+tmp[1033]*kernel[8];
				ans[933]<=tmp[832]*kernel[0]+tmp[833]*kernel[1]+tmp[834]*kernel[2]+tmp[932]*kernel[3]+tmp[933]*kernel[4]+tmp[934]*kernel[5]+tmp[1032]*kernel[6]+tmp[1033]*kernel[7]+tmp[1034]*kernel[8];
				ans[934]<=tmp[833]*kernel[0]+tmp[834]*kernel[1]+tmp[835]*kernel[2]+tmp[933]*kernel[3]+tmp[934]*kernel[4]+tmp[935]*kernel[5]+tmp[1033]*kernel[6]+tmp[1034]*kernel[7]+tmp[1035]*kernel[8];
				ans[935]<=tmp[834]*kernel[0]+tmp[835]*kernel[1]+tmp[836]*kernel[2]+tmp[934]*kernel[3]+tmp[935]*kernel[4]+tmp[936]*kernel[5]+tmp[1034]*kernel[6]+tmp[1035]*kernel[7]+tmp[1036]*kernel[8];
				ans[936]<=tmp[835]*kernel[0]+tmp[836]*kernel[1]+tmp[837]*kernel[2]+tmp[935]*kernel[3]+tmp[936]*kernel[4]+tmp[937]*kernel[5]+tmp[1035]*kernel[6]+tmp[1036]*kernel[7]+tmp[1037]*kernel[8];
				ans[937]<=tmp[836]*kernel[0]+tmp[837]*kernel[1]+tmp[838]*kernel[2]+tmp[936]*kernel[3]+tmp[937]*kernel[4]+tmp[938]*kernel[5]+tmp[1036]*kernel[6]+tmp[1037]*kernel[7]+tmp[1038]*kernel[8];
				ans[938]<=tmp[837]*kernel[0]+tmp[838]*kernel[1]+tmp[839]*kernel[2]+tmp[937]*kernel[3]+tmp[938]*kernel[4]+tmp[939]*kernel[5]+tmp[1037]*kernel[6]+tmp[1038]*kernel[7]+tmp[1039]*kernel[8];
				ans[939]<=tmp[838]*kernel[0]+tmp[839]*kernel[1]+tmp[840]*kernel[2]+tmp[938]*kernel[3]+tmp[939]*kernel[4]+tmp[940]*kernel[5]+tmp[1038]*kernel[6]+tmp[1039]*kernel[7]+tmp[1040]*kernel[8];
				ans[940]<=tmp[839]*kernel[0]+tmp[840]*kernel[1]+tmp[841]*kernel[2]+tmp[939]*kernel[3]+tmp[940]*kernel[4]+tmp[941]*kernel[5]+tmp[1039]*kernel[6]+tmp[1040]*kernel[7]+tmp[1041]*kernel[8];
				ans[941]<=tmp[840]*kernel[0]+tmp[841]*kernel[1]+tmp[842]*kernel[2]+tmp[940]*kernel[3]+tmp[941]*kernel[4]+tmp[942]*kernel[5]+tmp[1040]*kernel[6]+tmp[1041]*kernel[7]+tmp[1042]*kernel[8];
				ans[942]<=tmp[841]*kernel[0]+tmp[842]*kernel[1]+tmp[843]*kernel[2]+tmp[941]*kernel[3]+tmp[942]*kernel[4]+tmp[943]*kernel[5]+tmp[1041]*kernel[6]+tmp[1042]*kernel[7]+tmp[1043]*kernel[8];
				ans[943]<=tmp[842]*kernel[0]+tmp[843]*kernel[1]+tmp[844]*kernel[2]+tmp[942]*kernel[3]+tmp[943]*kernel[4]+tmp[944]*kernel[5]+tmp[1042]*kernel[6]+tmp[1043]*kernel[7]+tmp[1044]*kernel[8];
				ans[944]<=tmp[843]*kernel[0]+tmp[844]*kernel[1]+tmp[845]*kernel[2]+tmp[943]*kernel[3]+tmp[944]*kernel[4]+tmp[945]*kernel[5]+tmp[1043]*kernel[6]+tmp[1044]*kernel[7]+tmp[1045]*kernel[8];
				ans[945]<=tmp[844]*kernel[0]+tmp[845]*kernel[1]+tmp[846]*kernel[2]+tmp[944]*kernel[3]+tmp[945]*kernel[4]+tmp[946]*kernel[5]+tmp[1044]*kernel[6]+tmp[1045]*kernel[7]+tmp[1046]*kernel[8];
				ans[946]<=tmp[845]*kernel[0]+tmp[846]*kernel[1]+tmp[847]*kernel[2]+tmp[945]*kernel[3]+tmp[946]*kernel[4]+tmp[947]*kernel[5]+tmp[1045]*kernel[6]+tmp[1046]*kernel[7]+tmp[1047]*kernel[8];
				ans[947]<=tmp[846]*kernel[0]+tmp[847]*kernel[1]+tmp[848]*kernel[2]+tmp[946]*kernel[3]+tmp[947]*kernel[4]+tmp[948]*kernel[5]+tmp[1046]*kernel[6]+tmp[1047]*kernel[7]+tmp[1048]*kernel[8];
				ans[948]<=tmp[847]*kernel[0]+tmp[848]*kernel[1]+tmp[849]*kernel[2]+tmp[947]*kernel[3]+tmp[948]*kernel[4]+tmp[949]*kernel[5]+tmp[1047]*kernel[6]+tmp[1048]*kernel[7]+tmp[1049]*kernel[8];
				ans[949]<=tmp[848]*kernel[0]+tmp[849]*kernel[1]+tmp[850]*kernel[2]+tmp[948]*kernel[3]+tmp[949]*kernel[4]+tmp[950]*kernel[5]+tmp[1048]*kernel[6]+tmp[1049]*kernel[7]+tmp[1050]*kernel[8];
				ans[950]<=tmp[849]*kernel[0]+tmp[850]*kernel[1]+tmp[851]*kernel[2]+tmp[949]*kernel[3]+tmp[950]*kernel[4]+tmp[951]*kernel[5]+tmp[1049]*kernel[6]+tmp[1050]*kernel[7]+tmp[1051]*kernel[8];
				ans[951]<=tmp[850]*kernel[0]+tmp[851]*kernel[1]+tmp[852]*kernel[2]+tmp[950]*kernel[3]+tmp[951]*kernel[4]+tmp[952]*kernel[5]+tmp[1050]*kernel[6]+tmp[1051]*kernel[7]+tmp[1052]*kernel[8];
				ans[952]<=tmp[851]*kernel[0]+tmp[852]*kernel[1]+tmp[853]*kernel[2]+tmp[951]*kernel[3]+tmp[952]*kernel[4]+tmp[953]*kernel[5]+tmp[1051]*kernel[6]+tmp[1052]*kernel[7]+tmp[1053]*kernel[8];
				ans[953]<=tmp[852]*kernel[0]+tmp[853]*kernel[1]+tmp[854]*kernel[2]+tmp[952]*kernel[3]+tmp[953]*kernel[4]+tmp[954]*kernel[5]+tmp[1052]*kernel[6]+tmp[1053]*kernel[7]+tmp[1054]*kernel[8];
				ans[954]<=tmp[853]*kernel[0]+tmp[854]*kernel[1]+tmp[855]*kernel[2]+tmp[953]*kernel[3]+tmp[954]*kernel[4]+tmp[955]*kernel[5]+tmp[1053]*kernel[6]+tmp[1054]*kernel[7]+tmp[1055]*kernel[8];
				ans[955]<=tmp[854]*kernel[0]+tmp[855]*kernel[1]+tmp[856]*kernel[2]+tmp[954]*kernel[3]+tmp[955]*kernel[4]+tmp[956]*kernel[5]+tmp[1054]*kernel[6]+tmp[1055]*kernel[7]+tmp[1056]*kernel[8];
				ans[956]<=tmp[855]*kernel[0]+tmp[856]*kernel[1]+tmp[857]*kernel[2]+tmp[955]*kernel[3]+tmp[956]*kernel[4]+tmp[957]*kernel[5]+tmp[1055]*kernel[6]+tmp[1056]*kernel[7]+tmp[1057]*kernel[8];
				ans[957]<=tmp[856]*kernel[0]+tmp[857]*kernel[1]+tmp[858]*kernel[2]+tmp[956]*kernel[3]+tmp[957]*kernel[4]+tmp[958]*kernel[5]+tmp[1056]*kernel[6]+tmp[1057]*kernel[7]+tmp[1058]*kernel[8];
				ans[958]<=tmp[857]*kernel[0]+tmp[858]*kernel[1]+tmp[859]*kernel[2]+tmp[957]*kernel[3]+tmp[958]*kernel[4]+tmp[959]*kernel[5]+tmp[1057]*kernel[6]+tmp[1058]*kernel[7]+tmp[1059]*kernel[8];
				ans[959]<=tmp[858]*kernel[0]+tmp[859]*kernel[1]+tmp[860]*kernel[2]+tmp[958]*kernel[3]+tmp[959]*kernel[4]+tmp[960]*kernel[5]+tmp[1058]*kernel[6]+tmp[1059]*kernel[7]+tmp[1060]*kernel[8];
				ans[960]<=tmp[859]*kernel[0]+tmp[860]*kernel[1]+tmp[861]*kernel[2]+tmp[959]*kernel[3]+tmp[960]*kernel[4]+tmp[961]*kernel[5]+tmp[1059]*kernel[6]+tmp[1060]*kernel[7]+tmp[1061]*kernel[8];
				ans[961]<=tmp[860]*kernel[0]+tmp[861]*kernel[1]+tmp[862]*kernel[2]+tmp[960]*kernel[3]+tmp[961]*kernel[4]+tmp[962]*kernel[5]+tmp[1060]*kernel[6]+tmp[1061]*kernel[7]+tmp[1062]*kernel[8];
				ans[962]<=tmp[861]*kernel[0]+tmp[862]*kernel[1]+tmp[863]*kernel[2]+tmp[961]*kernel[3]+tmp[962]*kernel[4]+tmp[963]*kernel[5]+tmp[1061]*kernel[6]+tmp[1062]*kernel[7]+tmp[1063]*kernel[8];
				ans[963]<=tmp[862]*kernel[0]+tmp[863]*kernel[1]+tmp[864]*kernel[2]+tmp[962]*kernel[3]+tmp[963]*kernel[4]+tmp[964]*kernel[5]+tmp[1062]*kernel[6]+tmp[1063]*kernel[7]+tmp[1064]*kernel[8];
				ans[964]<=tmp[863]*kernel[0]+tmp[864]*kernel[1]+tmp[865]*kernel[2]+tmp[963]*kernel[3]+tmp[964]*kernel[4]+tmp[965]*kernel[5]+tmp[1063]*kernel[6]+tmp[1064]*kernel[7]+tmp[1065]*kernel[8];
				ans[965]<=tmp[864]*kernel[0]+tmp[865]*kernel[1]+tmp[866]*kernel[2]+tmp[964]*kernel[3]+tmp[965]*kernel[4]+tmp[966]*kernel[5]+tmp[1064]*kernel[6]+tmp[1065]*kernel[7]+tmp[1066]*kernel[8];
				ans[966]<=tmp[865]*kernel[0]+tmp[866]*kernel[1]+tmp[867]*kernel[2]+tmp[965]*kernel[3]+tmp[966]*kernel[4]+tmp[967]*kernel[5]+tmp[1065]*kernel[6]+tmp[1066]*kernel[7]+tmp[1067]*kernel[8];
				ans[967]<=tmp[866]*kernel[0]+tmp[867]*kernel[1]+tmp[868]*kernel[2]+tmp[966]*kernel[3]+tmp[967]*kernel[4]+tmp[968]*kernel[5]+tmp[1066]*kernel[6]+tmp[1067]*kernel[7]+tmp[1068]*kernel[8];
				ans[968]<=tmp[867]*kernel[0]+tmp[868]*kernel[1]+tmp[869]*kernel[2]+tmp[967]*kernel[3]+tmp[968]*kernel[4]+tmp[969]*kernel[5]+tmp[1067]*kernel[6]+tmp[1068]*kernel[7]+tmp[1069]*kernel[8];
				ans[969]<=tmp[868]*kernel[0]+tmp[869]*kernel[1]+tmp[870]*kernel[2]+tmp[968]*kernel[3]+tmp[969]*kernel[4]+tmp[970]*kernel[5]+tmp[1068]*kernel[6]+tmp[1069]*kernel[7]+tmp[1070]*kernel[8];
				ans[970]<=tmp[869]*kernel[0]+tmp[870]*kernel[1]+tmp[871]*kernel[2]+tmp[969]*kernel[3]+tmp[970]*kernel[4]+tmp[971]*kernel[5]+tmp[1069]*kernel[6]+tmp[1070]*kernel[7]+tmp[1071]*kernel[8];
				ans[971]<=tmp[870]*kernel[0]+tmp[871]*kernel[1]+tmp[872]*kernel[2]+tmp[970]*kernel[3]+tmp[971]*kernel[4]+tmp[972]*kernel[5]+tmp[1070]*kernel[6]+tmp[1071]*kernel[7]+tmp[1072]*kernel[8];
				ans[972]<=tmp[871]*kernel[0]+tmp[872]*kernel[1]+tmp[873]*kernel[2]+tmp[971]*kernel[3]+tmp[972]*kernel[4]+tmp[973]*kernel[5]+tmp[1071]*kernel[6]+tmp[1072]*kernel[7]+tmp[1073]*kernel[8];
				ans[973]<=tmp[872]*kernel[0]+tmp[873]*kernel[1]+tmp[874]*kernel[2]+tmp[972]*kernel[3]+tmp[973]*kernel[4]+tmp[974]*kernel[5]+tmp[1072]*kernel[6]+tmp[1073]*kernel[7]+tmp[1074]*kernel[8];
				ans[974]<=tmp[873]*kernel[0]+tmp[874]*kernel[1]+tmp[875]*kernel[2]+tmp[973]*kernel[3]+tmp[974]*kernel[4]+tmp[975]*kernel[5]+tmp[1073]*kernel[6]+tmp[1074]*kernel[7]+tmp[1075]*kernel[8];
				ans[975]<=tmp[874]*kernel[0]+tmp[875]*kernel[1]+tmp[876]*kernel[2]+tmp[974]*kernel[3]+tmp[975]*kernel[4]+tmp[976]*kernel[5]+tmp[1074]*kernel[6]+tmp[1075]*kernel[7]+tmp[1076]*kernel[8];
				ans[976]<=tmp[875]*kernel[0]+tmp[876]*kernel[1]+tmp[877]*kernel[2]+tmp[975]*kernel[3]+tmp[976]*kernel[4]+tmp[977]*kernel[5]+tmp[1075]*kernel[6]+tmp[1076]*kernel[7]+tmp[1077]*kernel[8];
				ans[977]<=tmp[876]*kernel[0]+tmp[877]*kernel[1]+tmp[878]*kernel[2]+tmp[976]*kernel[3]+tmp[977]*kernel[4]+tmp[978]*kernel[5]+tmp[1076]*kernel[6]+tmp[1077]*kernel[7]+tmp[1078]*kernel[8];
				ans[978]<=tmp[877]*kernel[0]+tmp[878]*kernel[1]+tmp[879]*kernel[2]+tmp[977]*kernel[3]+tmp[978]*kernel[4]+tmp[979]*kernel[5]+tmp[1077]*kernel[6]+tmp[1078]*kernel[7]+tmp[1079]*kernel[8];
				ans[979]<=tmp[878]*kernel[0]+tmp[879]*kernel[1]+tmp[880]*kernel[2]+tmp[978]*kernel[3]+tmp[979]*kernel[4]+tmp[980]*kernel[5]+tmp[1078]*kernel[6]+tmp[1079]*kernel[7]+tmp[1080]*kernel[8];
				ans[980]<=tmp[879]*kernel[0]+tmp[880]*kernel[1]+tmp[881]*kernel[2]+tmp[979]*kernel[3]+tmp[980]*kernel[4]+tmp[981]*kernel[5]+tmp[1079]*kernel[6]+tmp[1080]*kernel[7]+tmp[1081]*kernel[8];
				ans[981]<=tmp[880]*kernel[0]+tmp[881]*kernel[1]+tmp[882]*kernel[2]+tmp[980]*kernel[3]+tmp[981]*kernel[4]+tmp[982]*kernel[5]+tmp[1080]*kernel[6]+tmp[1081]*kernel[7]+tmp[1082]*kernel[8];
				ans[982]<=tmp[881]*kernel[0]+tmp[882]*kernel[1]+tmp[883]*kernel[2]+tmp[981]*kernel[3]+tmp[982]*kernel[4]+tmp[983]*kernel[5]+tmp[1081]*kernel[6]+tmp[1082]*kernel[7]+tmp[1083]*kernel[8];
				ans[983]<=tmp[882]*kernel[0]+tmp[883]*kernel[1]+tmp[884]*kernel[2]+tmp[982]*kernel[3]+tmp[983]*kernel[4]+tmp[984]*kernel[5]+tmp[1082]*kernel[6]+tmp[1083]*kernel[7]+tmp[1084]*kernel[8];
				ans[984]<=tmp[883]*kernel[0]+tmp[884]*kernel[1]+tmp[885]*kernel[2]+tmp[983]*kernel[3]+tmp[984]*kernel[4]+tmp[985]*kernel[5]+tmp[1083]*kernel[6]+tmp[1084]*kernel[7]+tmp[1085]*kernel[8];
				ans[985]<=tmp[884]*kernel[0]+tmp[885]*kernel[1]+tmp[886]*kernel[2]+tmp[984]*kernel[3]+tmp[985]*kernel[4]+tmp[986]*kernel[5]+tmp[1084]*kernel[6]+tmp[1085]*kernel[7]+tmp[1086]*kernel[8];
				ans[986]<=tmp[885]*kernel[0]+tmp[886]*kernel[1]+tmp[887]*kernel[2]+tmp[985]*kernel[3]+tmp[986]*kernel[4]+tmp[987]*kernel[5]+tmp[1085]*kernel[6]+tmp[1086]*kernel[7]+tmp[1087]*kernel[8];
				ans[987]<=tmp[886]*kernel[0]+tmp[887]*kernel[1]+tmp[888]*kernel[2]+tmp[986]*kernel[3]+tmp[987]*kernel[4]+tmp[988]*kernel[5]+tmp[1086]*kernel[6]+tmp[1087]*kernel[7]+tmp[1088]*kernel[8];
				ans[988]<=tmp[887]*kernel[0]+tmp[888]*kernel[1]+tmp[889]*kernel[2]+tmp[987]*kernel[3]+tmp[988]*kernel[4]+tmp[989]*kernel[5]+tmp[1087]*kernel[6]+tmp[1088]*kernel[7]+tmp[1089]*kernel[8];
				ans[989]<=tmp[888]*kernel[0]+tmp[889]*kernel[1]+tmp[890]*kernel[2]+tmp[988]*kernel[3]+tmp[989]*kernel[4]+tmp[990]*kernel[5]+tmp[1088]*kernel[6]+tmp[1089]*kernel[7]+tmp[1090]*kernel[8];
				ans[990]<=tmp[889]*kernel[0]+tmp[890]*kernel[1]+tmp[891]*kernel[2]+tmp[989]*kernel[3]+tmp[990]*kernel[4]+tmp[991]*kernel[5]+tmp[1089]*kernel[6]+tmp[1090]*kernel[7]+tmp[1091]*kernel[8];
				ans[991]<=tmp[890]*kernel[0]+tmp[891]*kernel[1]+tmp[892]*kernel[2]+tmp[990]*kernel[3]+tmp[991]*kernel[4]+tmp[992]*kernel[5]+tmp[1090]*kernel[6]+tmp[1091]*kernel[7]+tmp[1092]*kernel[8];
				ans[992]<=tmp[891]*kernel[0]+tmp[892]*kernel[1]+tmp[893]*kernel[2]+tmp[991]*kernel[3]+tmp[992]*kernel[4]+tmp[993]*kernel[5]+tmp[1091]*kernel[6]+tmp[1092]*kernel[7]+tmp[1093]*kernel[8];
				ans[993]<=tmp[892]*kernel[0]+tmp[893]*kernel[1]+tmp[894]*kernel[2]+tmp[992]*kernel[3]+tmp[993]*kernel[4]+tmp[994]*kernel[5]+tmp[1092]*kernel[6]+tmp[1093]*kernel[7]+tmp[1094]*kernel[8];
				ans[994]<=tmp[893]*kernel[0]+tmp[894]*kernel[1]+tmp[895]*kernel[2]+tmp[993]*kernel[3]+tmp[994]*kernel[4]+tmp[995]*kernel[5]+tmp[1093]*kernel[6]+tmp[1094]*kernel[7]+tmp[1095]*kernel[8];
				ans[995]<=tmp[894]*kernel[0]+tmp[895]*kernel[1]+tmp[896]*kernel[2]+tmp[994]*kernel[3]+tmp[995]*kernel[4]+tmp[996]*kernel[5]+tmp[1094]*kernel[6]+tmp[1095]*kernel[7]+tmp[1096]*kernel[8];
				ans[996]<=tmp[895]*kernel[0]+tmp[896]*kernel[1]+tmp[897]*kernel[2]+tmp[995]*kernel[3]+tmp[996]*kernel[4]+tmp[997]*kernel[5]+tmp[1095]*kernel[6]+tmp[1096]*kernel[7]+tmp[1097]*kernel[8];
				ans[997]<=tmp[896]*kernel[0]+tmp[897]*kernel[1]+tmp[898]*kernel[2]+tmp[996]*kernel[3]+tmp[997]*kernel[4]+tmp[998]*kernel[5]+tmp[1096]*kernel[6]+tmp[1097]*kernel[7]+tmp[1098]*kernel[8];
				ans[998]<=tmp[897]*kernel[0]+tmp[898]*kernel[1]+tmp[899]*kernel[2]+tmp[997]*kernel[3]+tmp[998]*kernel[4]+tmp[999]*kernel[5]+tmp[1097]*kernel[6]+tmp[1098]*kernel[7]+tmp[1099]*kernel[8];
				ans[999]<=tmp[898]*kernel[0]+tmp[899]*kernel[1]+tmp[998]*kernel[3]+tmp[999]*kernel[4]+tmp[1098]*kernel[6]+tmp[1099]*kernel[7];
				ans[1000]<=tmp[900]*kernel[1]+tmp[901]*kernel[2]+tmp[1000]*kernel[4]+tmp[1001]*kernel[5]+tmp[1100]*kernel[7]+tmp[1101]*kernel[8];
				ans[1001]<=tmp[900]*kernel[0]+tmp[901]*kernel[1]+tmp[902]*kernel[2]+tmp[1000]*kernel[3]+tmp[1001]*kernel[4]+tmp[1002]*kernel[5]+tmp[1100]*kernel[6]+tmp[1101]*kernel[7]+tmp[1102]*kernel[8];
				ans[1002]<=tmp[901]*kernel[0]+tmp[902]*kernel[1]+tmp[903]*kernel[2]+tmp[1001]*kernel[3]+tmp[1002]*kernel[4]+tmp[1003]*kernel[5]+tmp[1101]*kernel[6]+tmp[1102]*kernel[7]+tmp[1103]*kernel[8];
				ans[1003]<=tmp[902]*kernel[0]+tmp[903]*kernel[1]+tmp[904]*kernel[2]+tmp[1002]*kernel[3]+tmp[1003]*kernel[4]+tmp[1004]*kernel[5]+tmp[1102]*kernel[6]+tmp[1103]*kernel[7]+tmp[1104]*kernel[8];
				ans[1004]<=tmp[903]*kernel[0]+tmp[904]*kernel[1]+tmp[905]*kernel[2]+tmp[1003]*kernel[3]+tmp[1004]*kernel[4]+tmp[1005]*kernel[5]+tmp[1103]*kernel[6]+tmp[1104]*kernel[7]+tmp[1105]*kernel[8];
				ans[1005]<=tmp[904]*kernel[0]+tmp[905]*kernel[1]+tmp[906]*kernel[2]+tmp[1004]*kernel[3]+tmp[1005]*kernel[4]+tmp[1006]*kernel[5]+tmp[1104]*kernel[6]+tmp[1105]*kernel[7]+tmp[1106]*kernel[8];
				ans[1006]<=tmp[905]*kernel[0]+tmp[906]*kernel[1]+tmp[907]*kernel[2]+tmp[1005]*kernel[3]+tmp[1006]*kernel[4]+tmp[1007]*kernel[5]+tmp[1105]*kernel[6]+tmp[1106]*kernel[7]+tmp[1107]*kernel[8];
				ans[1007]<=tmp[906]*kernel[0]+tmp[907]*kernel[1]+tmp[908]*kernel[2]+tmp[1006]*kernel[3]+tmp[1007]*kernel[4]+tmp[1008]*kernel[5]+tmp[1106]*kernel[6]+tmp[1107]*kernel[7]+tmp[1108]*kernel[8];
				ans[1008]<=tmp[907]*kernel[0]+tmp[908]*kernel[1]+tmp[909]*kernel[2]+tmp[1007]*kernel[3]+tmp[1008]*kernel[4]+tmp[1009]*kernel[5]+tmp[1107]*kernel[6]+tmp[1108]*kernel[7]+tmp[1109]*kernel[8];
				ans[1009]<=tmp[908]*kernel[0]+tmp[909]*kernel[1]+tmp[910]*kernel[2]+tmp[1008]*kernel[3]+tmp[1009]*kernel[4]+tmp[1010]*kernel[5]+tmp[1108]*kernel[6]+tmp[1109]*kernel[7]+tmp[1110]*kernel[8];
				ans[1010]<=tmp[909]*kernel[0]+tmp[910]*kernel[1]+tmp[911]*kernel[2]+tmp[1009]*kernel[3]+tmp[1010]*kernel[4]+tmp[1011]*kernel[5]+tmp[1109]*kernel[6]+tmp[1110]*kernel[7]+tmp[1111]*kernel[8];
				ans[1011]<=tmp[910]*kernel[0]+tmp[911]*kernel[1]+tmp[912]*kernel[2]+tmp[1010]*kernel[3]+tmp[1011]*kernel[4]+tmp[1012]*kernel[5]+tmp[1110]*kernel[6]+tmp[1111]*kernel[7]+tmp[1112]*kernel[8];
				ans[1012]<=tmp[911]*kernel[0]+tmp[912]*kernel[1]+tmp[913]*kernel[2]+tmp[1011]*kernel[3]+tmp[1012]*kernel[4]+tmp[1013]*kernel[5]+tmp[1111]*kernel[6]+tmp[1112]*kernel[7]+tmp[1113]*kernel[8];
				ans[1013]<=tmp[912]*kernel[0]+tmp[913]*kernel[1]+tmp[914]*kernel[2]+tmp[1012]*kernel[3]+tmp[1013]*kernel[4]+tmp[1014]*kernel[5]+tmp[1112]*kernel[6]+tmp[1113]*kernel[7]+tmp[1114]*kernel[8];
				ans[1014]<=tmp[913]*kernel[0]+tmp[914]*kernel[1]+tmp[915]*kernel[2]+tmp[1013]*kernel[3]+tmp[1014]*kernel[4]+tmp[1015]*kernel[5]+tmp[1113]*kernel[6]+tmp[1114]*kernel[7]+tmp[1115]*kernel[8];
				ans[1015]<=tmp[914]*kernel[0]+tmp[915]*kernel[1]+tmp[916]*kernel[2]+tmp[1014]*kernel[3]+tmp[1015]*kernel[4]+tmp[1016]*kernel[5]+tmp[1114]*kernel[6]+tmp[1115]*kernel[7]+tmp[1116]*kernel[8];
				ans[1016]<=tmp[915]*kernel[0]+tmp[916]*kernel[1]+tmp[917]*kernel[2]+tmp[1015]*kernel[3]+tmp[1016]*kernel[4]+tmp[1017]*kernel[5]+tmp[1115]*kernel[6]+tmp[1116]*kernel[7]+tmp[1117]*kernel[8];
				ans[1017]<=tmp[916]*kernel[0]+tmp[917]*kernel[1]+tmp[918]*kernel[2]+tmp[1016]*kernel[3]+tmp[1017]*kernel[4]+tmp[1018]*kernel[5]+tmp[1116]*kernel[6]+tmp[1117]*kernel[7]+tmp[1118]*kernel[8];
				ans[1018]<=tmp[917]*kernel[0]+tmp[918]*kernel[1]+tmp[919]*kernel[2]+tmp[1017]*kernel[3]+tmp[1018]*kernel[4]+tmp[1019]*kernel[5]+tmp[1117]*kernel[6]+tmp[1118]*kernel[7]+tmp[1119]*kernel[8];
				ans[1019]<=tmp[918]*kernel[0]+tmp[919]*kernel[1]+tmp[920]*kernel[2]+tmp[1018]*kernel[3]+tmp[1019]*kernel[4]+tmp[1020]*kernel[5]+tmp[1118]*kernel[6]+tmp[1119]*kernel[7]+tmp[1120]*kernel[8];
				ans[1020]<=tmp[919]*kernel[0]+tmp[920]*kernel[1]+tmp[921]*kernel[2]+tmp[1019]*kernel[3]+tmp[1020]*kernel[4]+tmp[1021]*kernel[5]+tmp[1119]*kernel[6]+tmp[1120]*kernel[7]+tmp[1121]*kernel[8];
				ans[1021]<=tmp[920]*kernel[0]+tmp[921]*kernel[1]+tmp[922]*kernel[2]+tmp[1020]*kernel[3]+tmp[1021]*kernel[4]+tmp[1022]*kernel[5]+tmp[1120]*kernel[6]+tmp[1121]*kernel[7]+tmp[1122]*kernel[8];
				ans[1022]<=tmp[921]*kernel[0]+tmp[922]*kernel[1]+tmp[923]*kernel[2]+tmp[1021]*kernel[3]+tmp[1022]*kernel[4]+tmp[1023]*kernel[5]+tmp[1121]*kernel[6]+tmp[1122]*kernel[7]+tmp[1123]*kernel[8];
				ans[1023]<=tmp[922]*kernel[0]+tmp[923]*kernel[1]+tmp[924]*kernel[2]+tmp[1022]*kernel[3]+tmp[1023]*kernel[4]+tmp[1024]*kernel[5]+tmp[1122]*kernel[6]+tmp[1123]*kernel[7]+tmp[1124]*kernel[8];
				ans[1024]<=tmp[923]*kernel[0]+tmp[924]*kernel[1]+tmp[925]*kernel[2]+tmp[1023]*kernel[3]+tmp[1024]*kernel[4]+tmp[1025]*kernel[5]+tmp[1123]*kernel[6]+tmp[1124]*kernel[7]+tmp[1125]*kernel[8];
				ans[1025]<=tmp[924]*kernel[0]+tmp[925]*kernel[1]+tmp[926]*kernel[2]+tmp[1024]*kernel[3]+tmp[1025]*kernel[4]+tmp[1026]*kernel[5]+tmp[1124]*kernel[6]+tmp[1125]*kernel[7]+tmp[1126]*kernel[8];
				ans[1026]<=tmp[925]*kernel[0]+tmp[926]*kernel[1]+tmp[927]*kernel[2]+tmp[1025]*kernel[3]+tmp[1026]*kernel[4]+tmp[1027]*kernel[5]+tmp[1125]*kernel[6]+tmp[1126]*kernel[7]+tmp[1127]*kernel[8];
				ans[1027]<=tmp[926]*kernel[0]+tmp[927]*kernel[1]+tmp[928]*kernel[2]+tmp[1026]*kernel[3]+tmp[1027]*kernel[4]+tmp[1028]*kernel[5]+tmp[1126]*kernel[6]+tmp[1127]*kernel[7]+tmp[1128]*kernel[8];
				ans[1028]<=tmp[927]*kernel[0]+tmp[928]*kernel[1]+tmp[929]*kernel[2]+tmp[1027]*kernel[3]+tmp[1028]*kernel[4]+tmp[1029]*kernel[5]+tmp[1127]*kernel[6]+tmp[1128]*kernel[7]+tmp[1129]*kernel[8];
				ans[1029]<=tmp[928]*kernel[0]+tmp[929]*kernel[1]+tmp[930]*kernel[2]+tmp[1028]*kernel[3]+tmp[1029]*kernel[4]+tmp[1030]*kernel[5]+tmp[1128]*kernel[6]+tmp[1129]*kernel[7]+tmp[1130]*kernel[8];
				ans[1030]<=tmp[929]*kernel[0]+tmp[930]*kernel[1]+tmp[931]*kernel[2]+tmp[1029]*kernel[3]+tmp[1030]*kernel[4]+tmp[1031]*kernel[5]+tmp[1129]*kernel[6]+tmp[1130]*kernel[7]+tmp[1131]*kernel[8];
				ans[1031]<=tmp[930]*kernel[0]+tmp[931]*kernel[1]+tmp[932]*kernel[2]+tmp[1030]*kernel[3]+tmp[1031]*kernel[4]+tmp[1032]*kernel[5]+tmp[1130]*kernel[6]+tmp[1131]*kernel[7]+tmp[1132]*kernel[8];
				ans[1032]<=tmp[931]*kernel[0]+tmp[932]*kernel[1]+tmp[933]*kernel[2]+tmp[1031]*kernel[3]+tmp[1032]*kernel[4]+tmp[1033]*kernel[5]+tmp[1131]*kernel[6]+tmp[1132]*kernel[7]+tmp[1133]*kernel[8];
				ans[1033]<=tmp[932]*kernel[0]+tmp[933]*kernel[1]+tmp[934]*kernel[2]+tmp[1032]*kernel[3]+tmp[1033]*kernel[4]+tmp[1034]*kernel[5]+tmp[1132]*kernel[6]+tmp[1133]*kernel[7]+tmp[1134]*kernel[8];
				ans[1034]<=tmp[933]*kernel[0]+tmp[934]*kernel[1]+tmp[935]*kernel[2]+tmp[1033]*kernel[3]+tmp[1034]*kernel[4]+tmp[1035]*kernel[5]+tmp[1133]*kernel[6]+tmp[1134]*kernel[7]+tmp[1135]*kernel[8];
				ans[1035]<=tmp[934]*kernel[0]+tmp[935]*kernel[1]+tmp[936]*kernel[2]+tmp[1034]*kernel[3]+tmp[1035]*kernel[4]+tmp[1036]*kernel[5]+tmp[1134]*kernel[6]+tmp[1135]*kernel[7]+tmp[1136]*kernel[8];
				ans[1036]<=tmp[935]*kernel[0]+tmp[936]*kernel[1]+tmp[937]*kernel[2]+tmp[1035]*kernel[3]+tmp[1036]*kernel[4]+tmp[1037]*kernel[5]+tmp[1135]*kernel[6]+tmp[1136]*kernel[7]+tmp[1137]*kernel[8];
				ans[1037]<=tmp[936]*kernel[0]+tmp[937]*kernel[1]+tmp[938]*kernel[2]+tmp[1036]*kernel[3]+tmp[1037]*kernel[4]+tmp[1038]*kernel[5]+tmp[1136]*kernel[6]+tmp[1137]*kernel[7]+tmp[1138]*kernel[8];
				ans[1038]<=tmp[937]*kernel[0]+tmp[938]*kernel[1]+tmp[939]*kernel[2]+tmp[1037]*kernel[3]+tmp[1038]*kernel[4]+tmp[1039]*kernel[5]+tmp[1137]*kernel[6]+tmp[1138]*kernel[7]+tmp[1139]*kernel[8];
				ans[1039]<=tmp[938]*kernel[0]+tmp[939]*kernel[1]+tmp[940]*kernel[2]+tmp[1038]*kernel[3]+tmp[1039]*kernel[4]+tmp[1040]*kernel[5]+tmp[1138]*kernel[6]+tmp[1139]*kernel[7]+tmp[1140]*kernel[8];
				ans[1040]<=tmp[939]*kernel[0]+tmp[940]*kernel[1]+tmp[941]*kernel[2]+tmp[1039]*kernel[3]+tmp[1040]*kernel[4]+tmp[1041]*kernel[5]+tmp[1139]*kernel[6]+tmp[1140]*kernel[7]+tmp[1141]*kernel[8];
				ans[1041]<=tmp[940]*kernel[0]+tmp[941]*kernel[1]+tmp[942]*kernel[2]+tmp[1040]*kernel[3]+tmp[1041]*kernel[4]+tmp[1042]*kernel[5]+tmp[1140]*kernel[6]+tmp[1141]*kernel[7]+tmp[1142]*kernel[8];
				ans[1042]<=tmp[941]*kernel[0]+tmp[942]*kernel[1]+tmp[943]*kernel[2]+tmp[1041]*kernel[3]+tmp[1042]*kernel[4]+tmp[1043]*kernel[5]+tmp[1141]*kernel[6]+tmp[1142]*kernel[7]+tmp[1143]*kernel[8];
				ans[1043]<=tmp[942]*kernel[0]+tmp[943]*kernel[1]+tmp[944]*kernel[2]+tmp[1042]*kernel[3]+tmp[1043]*kernel[4]+tmp[1044]*kernel[5]+tmp[1142]*kernel[6]+tmp[1143]*kernel[7]+tmp[1144]*kernel[8];
				ans[1044]<=tmp[943]*kernel[0]+tmp[944]*kernel[1]+tmp[945]*kernel[2]+tmp[1043]*kernel[3]+tmp[1044]*kernel[4]+tmp[1045]*kernel[5]+tmp[1143]*kernel[6]+tmp[1144]*kernel[7]+tmp[1145]*kernel[8];
				ans[1045]<=tmp[944]*kernel[0]+tmp[945]*kernel[1]+tmp[946]*kernel[2]+tmp[1044]*kernel[3]+tmp[1045]*kernel[4]+tmp[1046]*kernel[5]+tmp[1144]*kernel[6]+tmp[1145]*kernel[7]+tmp[1146]*kernel[8];
				ans[1046]<=tmp[945]*kernel[0]+tmp[946]*kernel[1]+tmp[947]*kernel[2]+tmp[1045]*kernel[3]+tmp[1046]*kernel[4]+tmp[1047]*kernel[5]+tmp[1145]*kernel[6]+tmp[1146]*kernel[7]+tmp[1147]*kernel[8];
				ans[1047]<=tmp[946]*kernel[0]+tmp[947]*kernel[1]+tmp[948]*kernel[2]+tmp[1046]*kernel[3]+tmp[1047]*kernel[4]+tmp[1048]*kernel[5]+tmp[1146]*kernel[6]+tmp[1147]*kernel[7]+tmp[1148]*kernel[8];
				ans[1048]<=tmp[947]*kernel[0]+tmp[948]*kernel[1]+tmp[949]*kernel[2]+tmp[1047]*kernel[3]+tmp[1048]*kernel[4]+tmp[1049]*kernel[5]+tmp[1147]*kernel[6]+tmp[1148]*kernel[7]+tmp[1149]*kernel[8];
				ans[1049]<=tmp[948]*kernel[0]+tmp[949]*kernel[1]+tmp[950]*kernel[2]+tmp[1048]*kernel[3]+tmp[1049]*kernel[4]+tmp[1050]*kernel[5]+tmp[1148]*kernel[6]+tmp[1149]*kernel[7]+tmp[1150]*kernel[8];
				ans[1050]<=tmp[949]*kernel[0]+tmp[950]*kernel[1]+tmp[951]*kernel[2]+tmp[1049]*kernel[3]+tmp[1050]*kernel[4]+tmp[1051]*kernel[5]+tmp[1149]*kernel[6]+tmp[1150]*kernel[7]+tmp[1151]*kernel[8];
				ans[1051]<=tmp[950]*kernel[0]+tmp[951]*kernel[1]+tmp[952]*kernel[2]+tmp[1050]*kernel[3]+tmp[1051]*kernel[4]+tmp[1052]*kernel[5]+tmp[1150]*kernel[6]+tmp[1151]*kernel[7]+tmp[1152]*kernel[8];
				ans[1052]<=tmp[951]*kernel[0]+tmp[952]*kernel[1]+tmp[953]*kernel[2]+tmp[1051]*kernel[3]+tmp[1052]*kernel[4]+tmp[1053]*kernel[5]+tmp[1151]*kernel[6]+tmp[1152]*kernel[7]+tmp[1153]*kernel[8];
				ans[1053]<=tmp[952]*kernel[0]+tmp[953]*kernel[1]+tmp[954]*kernel[2]+tmp[1052]*kernel[3]+tmp[1053]*kernel[4]+tmp[1054]*kernel[5]+tmp[1152]*kernel[6]+tmp[1153]*kernel[7]+tmp[1154]*kernel[8];
				ans[1054]<=tmp[953]*kernel[0]+tmp[954]*kernel[1]+tmp[955]*kernel[2]+tmp[1053]*kernel[3]+tmp[1054]*kernel[4]+tmp[1055]*kernel[5]+tmp[1153]*kernel[6]+tmp[1154]*kernel[7]+tmp[1155]*kernel[8];
				ans[1055]<=tmp[954]*kernel[0]+tmp[955]*kernel[1]+tmp[956]*kernel[2]+tmp[1054]*kernel[3]+tmp[1055]*kernel[4]+tmp[1056]*kernel[5]+tmp[1154]*kernel[6]+tmp[1155]*kernel[7]+tmp[1156]*kernel[8];
				ans[1056]<=tmp[955]*kernel[0]+tmp[956]*kernel[1]+tmp[957]*kernel[2]+tmp[1055]*kernel[3]+tmp[1056]*kernel[4]+tmp[1057]*kernel[5]+tmp[1155]*kernel[6]+tmp[1156]*kernel[7]+tmp[1157]*kernel[8];
				ans[1057]<=tmp[956]*kernel[0]+tmp[957]*kernel[1]+tmp[958]*kernel[2]+tmp[1056]*kernel[3]+tmp[1057]*kernel[4]+tmp[1058]*kernel[5]+tmp[1156]*kernel[6]+tmp[1157]*kernel[7]+tmp[1158]*kernel[8];
				ans[1058]<=tmp[957]*kernel[0]+tmp[958]*kernel[1]+tmp[959]*kernel[2]+tmp[1057]*kernel[3]+tmp[1058]*kernel[4]+tmp[1059]*kernel[5]+tmp[1157]*kernel[6]+tmp[1158]*kernel[7]+tmp[1159]*kernel[8];
				ans[1059]<=tmp[958]*kernel[0]+tmp[959]*kernel[1]+tmp[960]*kernel[2]+tmp[1058]*kernel[3]+tmp[1059]*kernel[4]+tmp[1060]*kernel[5]+tmp[1158]*kernel[6]+tmp[1159]*kernel[7]+tmp[1160]*kernel[8];
				ans[1060]<=tmp[959]*kernel[0]+tmp[960]*kernel[1]+tmp[961]*kernel[2]+tmp[1059]*kernel[3]+tmp[1060]*kernel[4]+tmp[1061]*kernel[5]+tmp[1159]*kernel[6]+tmp[1160]*kernel[7]+tmp[1161]*kernel[8];
				ans[1061]<=tmp[960]*kernel[0]+tmp[961]*kernel[1]+tmp[962]*kernel[2]+tmp[1060]*kernel[3]+tmp[1061]*kernel[4]+tmp[1062]*kernel[5]+tmp[1160]*kernel[6]+tmp[1161]*kernel[7]+tmp[1162]*kernel[8];
				ans[1062]<=tmp[961]*kernel[0]+tmp[962]*kernel[1]+tmp[963]*kernel[2]+tmp[1061]*kernel[3]+tmp[1062]*kernel[4]+tmp[1063]*kernel[5]+tmp[1161]*kernel[6]+tmp[1162]*kernel[7]+tmp[1163]*kernel[8];
				ans[1063]<=tmp[962]*kernel[0]+tmp[963]*kernel[1]+tmp[964]*kernel[2]+tmp[1062]*kernel[3]+tmp[1063]*kernel[4]+tmp[1064]*kernel[5]+tmp[1162]*kernel[6]+tmp[1163]*kernel[7]+tmp[1164]*kernel[8];
				ans[1064]<=tmp[963]*kernel[0]+tmp[964]*kernel[1]+tmp[965]*kernel[2]+tmp[1063]*kernel[3]+tmp[1064]*kernel[4]+tmp[1065]*kernel[5]+tmp[1163]*kernel[6]+tmp[1164]*kernel[7]+tmp[1165]*kernel[8];
				ans[1065]<=tmp[964]*kernel[0]+tmp[965]*kernel[1]+tmp[966]*kernel[2]+tmp[1064]*kernel[3]+tmp[1065]*kernel[4]+tmp[1066]*kernel[5]+tmp[1164]*kernel[6]+tmp[1165]*kernel[7]+tmp[1166]*kernel[8];
				ans[1066]<=tmp[965]*kernel[0]+tmp[966]*kernel[1]+tmp[967]*kernel[2]+tmp[1065]*kernel[3]+tmp[1066]*kernel[4]+tmp[1067]*kernel[5]+tmp[1165]*kernel[6]+tmp[1166]*kernel[7]+tmp[1167]*kernel[8];
				ans[1067]<=tmp[966]*kernel[0]+tmp[967]*kernel[1]+tmp[968]*kernel[2]+tmp[1066]*kernel[3]+tmp[1067]*kernel[4]+tmp[1068]*kernel[5]+tmp[1166]*kernel[6]+tmp[1167]*kernel[7]+tmp[1168]*kernel[8];
				ans[1068]<=tmp[967]*kernel[0]+tmp[968]*kernel[1]+tmp[969]*kernel[2]+tmp[1067]*kernel[3]+tmp[1068]*kernel[4]+tmp[1069]*kernel[5]+tmp[1167]*kernel[6]+tmp[1168]*kernel[7]+tmp[1169]*kernel[8];
				ans[1069]<=tmp[968]*kernel[0]+tmp[969]*kernel[1]+tmp[970]*kernel[2]+tmp[1068]*kernel[3]+tmp[1069]*kernel[4]+tmp[1070]*kernel[5]+tmp[1168]*kernel[6]+tmp[1169]*kernel[7]+tmp[1170]*kernel[8];
				ans[1070]<=tmp[969]*kernel[0]+tmp[970]*kernel[1]+tmp[971]*kernel[2]+tmp[1069]*kernel[3]+tmp[1070]*kernel[4]+tmp[1071]*kernel[5]+tmp[1169]*kernel[6]+tmp[1170]*kernel[7]+tmp[1171]*kernel[8];
				ans[1071]<=tmp[970]*kernel[0]+tmp[971]*kernel[1]+tmp[972]*kernel[2]+tmp[1070]*kernel[3]+tmp[1071]*kernel[4]+tmp[1072]*kernel[5]+tmp[1170]*kernel[6]+tmp[1171]*kernel[7]+tmp[1172]*kernel[8];
				ans[1072]<=tmp[971]*kernel[0]+tmp[972]*kernel[1]+tmp[973]*kernel[2]+tmp[1071]*kernel[3]+tmp[1072]*kernel[4]+tmp[1073]*kernel[5]+tmp[1171]*kernel[6]+tmp[1172]*kernel[7]+tmp[1173]*kernel[8];
				ans[1073]<=tmp[972]*kernel[0]+tmp[973]*kernel[1]+tmp[974]*kernel[2]+tmp[1072]*kernel[3]+tmp[1073]*kernel[4]+tmp[1074]*kernel[5]+tmp[1172]*kernel[6]+tmp[1173]*kernel[7]+tmp[1174]*kernel[8];
				ans[1074]<=tmp[973]*kernel[0]+tmp[974]*kernel[1]+tmp[975]*kernel[2]+tmp[1073]*kernel[3]+tmp[1074]*kernel[4]+tmp[1075]*kernel[5]+tmp[1173]*kernel[6]+tmp[1174]*kernel[7]+tmp[1175]*kernel[8];
				ans[1075]<=tmp[974]*kernel[0]+tmp[975]*kernel[1]+tmp[976]*kernel[2]+tmp[1074]*kernel[3]+tmp[1075]*kernel[4]+tmp[1076]*kernel[5]+tmp[1174]*kernel[6]+tmp[1175]*kernel[7]+tmp[1176]*kernel[8];
				ans[1076]<=tmp[975]*kernel[0]+tmp[976]*kernel[1]+tmp[977]*kernel[2]+tmp[1075]*kernel[3]+tmp[1076]*kernel[4]+tmp[1077]*kernel[5]+tmp[1175]*kernel[6]+tmp[1176]*kernel[7]+tmp[1177]*kernel[8];
				ans[1077]<=tmp[976]*kernel[0]+tmp[977]*kernel[1]+tmp[978]*kernel[2]+tmp[1076]*kernel[3]+tmp[1077]*kernel[4]+tmp[1078]*kernel[5]+tmp[1176]*kernel[6]+tmp[1177]*kernel[7]+tmp[1178]*kernel[8];
				ans[1078]<=tmp[977]*kernel[0]+tmp[978]*kernel[1]+tmp[979]*kernel[2]+tmp[1077]*kernel[3]+tmp[1078]*kernel[4]+tmp[1079]*kernel[5]+tmp[1177]*kernel[6]+tmp[1178]*kernel[7]+tmp[1179]*kernel[8];
				ans[1079]<=tmp[978]*kernel[0]+tmp[979]*kernel[1]+tmp[980]*kernel[2]+tmp[1078]*kernel[3]+tmp[1079]*kernel[4]+tmp[1080]*kernel[5]+tmp[1178]*kernel[6]+tmp[1179]*kernel[7]+tmp[1180]*kernel[8];
				ans[1080]<=tmp[979]*kernel[0]+tmp[980]*kernel[1]+tmp[981]*kernel[2]+tmp[1079]*kernel[3]+tmp[1080]*kernel[4]+tmp[1081]*kernel[5]+tmp[1179]*kernel[6]+tmp[1180]*kernel[7]+tmp[1181]*kernel[8];
				ans[1081]<=tmp[980]*kernel[0]+tmp[981]*kernel[1]+tmp[982]*kernel[2]+tmp[1080]*kernel[3]+tmp[1081]*kernel[4]+tmp[1082]*kernel[5]+tmp[1180]*kernel[6]+tmp[1181]*kernel[7]+tmp[1182]*kernel[8];
				ans[1082]<=tmp[981]*kernel[0]+tmp[982]*kernel[1]+tmp[983]*kernel[2]+tmp[1081]*kernel[3]+tmp[1082]*kernel[4]+tmp[1083]*kernel[5]+tmp[1181]*kernel[6]+tmp[1182]*kernel[7]+tmp[1183]*kernel[8];
				ans[1083]<=tmp[982]*kernel[0]+tmp[983]*kernel[1]+tmp[984]*kernel[2]+tmp[1082]*kernel[3]+tmp[1083]*kernel[4]+tmp[1084]*kernel[5]+tmp[1182]*kernel[6]+tmp[1183]*kernel[7]+tmp[1184]*kernel[8];
				ans[1084]<=tmp[983]*kernel[0]+tmp[984]*kernel[1]+tmp[985]*kernel[2]+tmp[1083]*kernel[3]+tmp[1084]*kernel[4]+tmp[1085]*kernel[5]+tmp[1183]*kernel[6]+tmp[1184]*kernel[7]+tmp[1185]*kernel[8];
				ans[1085]<=tmp[984]*kernel[0]+tmp[985]*kernel[1]+tmp[986]*kernel[2]+tmp[1084]*kernel[3]+tmp[1085]*kernel[4]+tmp[1086]*kernel[5]+tmp[1184]*kernel[6]+tmp[1185]*kernel[7]+tmp[1186]*kernel[8];
				ans[1086]<=tmp[985]*kernel[0]+tmp[986]*kernel[1]+tmp[987]*kernel[2]+tmp[1085]*kernel[3]+tmp[1086]*kernel[4]+tmp[1087]*kernel[5]+tmp[1185]*kernel[6]+tmp[1186]*kernel[7]+tmp[1187]*kernel[8];
				ans[1087]<=tmp[986]*kernel[0]+tmp[987]*kernel[1]+tmp[988]*kernel[2]+tmp[1086]*kernel[3]+tmp[1087]*kernel[4]+tmp[1088]*kernel[5]+tmp[1186]*kernel[6]+tmp[1187]*kernel[7]+tmp[1188]*kernel[8];
				ans[1088]<=tmp[987]*kernel[0]+tmp[988]*kernel[1]+tmp[989]*kernel[2]+tmp[1087]*kernel[3]+tmp[1088]*kernel[4]+tmp[1089]*kernel[5]+tmp[1187]*kernel[6]+tmp[1188]*kernel[7]+tmp[1189]*kernel[8];
				ans[1089]<=tmp[988]*kernel[0]+tmp[989]*kernel[1]+tmp[990]*kernel[2]+tmp[1088]*kernel[3]+tmp[1089]*kernel[4]+tmp[1090]*kernel[5]+tmp[1188]*kernel[6]+tmp[1189]*kernel[7]+tmp[1190]*kernel[8];
				ans[1090]<=tmp[989]*kernel[0]+tmp[990]*kernel[1]+tmp[991]*kernel[2]+tmp[1089]*kernel[3]+tmp[1090]*kernel[4]+tmp[1091]*kernel[5]+tmp[1189]*kernel[6]+tmp[1190]*kernel[7]+tmp[1191]*kernel[8];
				ans[1091]<=tmp[990]*kernel[0]+tmp[991]*kernel[1]+tmp[992]*kernel[2]+tmp[1090]*kernel[3]+tmp[1091]*kernel[4]+tmp[1092]*kernel[5]+tmp[1190]*kernel[6]+tmp[1191]*kernel[7]+tmp[1192]*kernel[8];
				ans[1092]<=tmp[991]*kernel[0]+tmp[992]*kernel[1]+tmp[993]*kernel[2]+tmp[1091]*kernel[3]+tmp[1092]*kernel[4]+tmp[1093]*kernel[5]+tmp[1191]*kernel[6]+tmp[1192]*kernel[7]+tmp[1193]*kernel[8];
				ans[1093]<=tmp[992]*kernel[0]+tmp[993]*kernel[1]+tmp[994]*kernel[2]+tmp[1092]*kernel[3]+tmp[1093]*kernel[4]+tmp[1094]*kernel[5]+tmp[1192]*kernel[6]+tmp[1193]*kernel[7]+tmp[1194]*kernel[8];
				ans[1094]<=tmp[993]*kernel[0]+tmp[994]*kernel[1]+tmp[995]*kernel[2]+tmp[1093]*kernel[3]+tmp[1094]*kernel[4]+tmp[1095]*kernel[5]+tmp[1193]*kernel[6]+tmp[1194]*kernel[7]+tmp[1195]*kernel[8];
				ans[1095]<=tmp[994]*kernel[0]+tmp[995]*kernel[1]+tmp[996]*kernel[2]+tmp[1094]*kernel[3]+tmp[1095]*kernel[4]+tmp[1096]*kernel[5]+tmp[1194]*kernel[6]+tmp[1195]*kernel[7]+tmp[1196]*kernel[8];
				ans[1096]<=tmp[995]*kernel[0]+tmp[996]*kernel[1]+tmp[997]*kernel[2]+tmp[1095]*kernel[3]+tmp[1096]*kernel[4]+tmp[1097]*kernel[5]+tmp[1195]*kernel[6]+tmp[1196]*kernel[7]+tmp[1197]*kernel[8];
				ans[1097]<=tmp[996]*kernel[0]+tmp[997]*kernel[1]+tmp[998]*kernel[2]+tmp[1096]*kernel[3]+tmp[1097]*kernel[4]+tmp[1098]*kernel[5]+tmp[1196]*kernel[6]+tmp[1197]*kernel[7]+tmp[1198]*kernel[8];
				ans[1098]<=tmp[997]*kernel[0]+tmp[998]*kernel[1]+tmp[999]*kernel[2]+tmp[1097]*kernel[3]+tmp[1098]*kernel[4]+tmp[1099]*kernel[5]+tmp[1197]*kernel[6]+tmp[1198]*kernel[7]+tmp[1199]*kernel[8];
				ans[1099]<=tmp[998]*kernel[0]+tmp[999]*kernel[1]+tmp[1098]*kernel[3]+tmp[1099]*kernel[4]+tmp[1198]*kernel[6]+tmp[1199]*kernel[7];
				ans[1100]<=tmp[1000]*kernel[1]+tmp[1001]*kernel[2]+tmp[1100]*kernel[4]+tmp[1101]*kernel[5]+tmp[1200]*kernel[7]+tmp[1201]*kernel[8];
				ans[1101]<=tmp[1000]*kernel[0]+tmp[1001]*kernel[1]+tmp[1002]*kernel[2]+tmp[1100]*kernel[3]+tmp[1101]*kernel[4]+tmp[1102]*kernel[5]+tmp[1200]*kernel[6]+tmp[1201]*kernel[7]+tmp[1202]*kernel[8];
				ans[1102]<=tmp[1001]*kernel[0]+tmp[1002]*kernel[1]+tmp[1003]*kernel[2]+tmp[1101]*kernel[3]+tmp[1102]*kernel[4]+tmp[1103]*kernel[5]+tmp[1201]*kernel[6]+tmp[1202]*kernel[7]+tmp[1203]*kernel[8];
				ans[1103]<=tmp[1002]*kernel[0]+tmp[1003]*kernel[1]+tmp[1004]*kernel[2]+tmp[1102]*kernel[3]+tmp[1103]*kernel[4]+tmp[1104]*kernel[5]+tmp[1202]*kernel[6]+tmp[1203]*kernel[7]+tmp[1204]*kernel[8];
				ans[1104]<=tmp[1003]*kernel[0]+tmp[1004]*kernel[1]+tmp[1005]*kernel[2]+tmp[1103]*kernel[3]+tmp[1104]*kernel[4]+tmp[1105]*kernel[5]+tmp[1203]*kernel[6]+tmp[1204]*kernel[7]+tmp[1205]*kernel[8];
				ans[1105]<=tmp[1004]*kernel[0]+tmp[1005]*kernel[1]+tmp[1006]*kernel[2]+tmp[1104]*kernel[3]+tmp[1105]*kernel[4]+tmp[1106]*kernel[5]+tmp[1204]*kernel[6]+tmp[1205]*kernel[7]+tmp[1206]*kernel[8];
				ans[1106]<=tmp[1005]*kernel[0]+tmp[1006]*kernel[1]+tmp[1007]*kernel[2]+tmp[1105]*kernel[3]+tmp[1106]*kernel[4]+tmp[1107]*kernel[5]+tmp[1205]*kernel[6]+tmp[1206]*kernel[7]+tmp[1207]*kernel[8];
				ans[1107]<=tmp[1006]*kernel[0]+tmp[1007]*kernel[1]+tmp[1008]*kernel[2]+tmp[1106]*kernel[3]+tmp[1107]*kernel[4]+tmp[1108]*kernel[5]+tmp[1206]*kernel[6]+tmp[1207]*kernel[7]+tmp[1208]*kernel[8];
				ans[1108]<=tmp[1007]*kernel[0]+tmp[1008]*kernel[1]+tmp[1009]*kernel[2]+tmp[1107]*kernel[3]+tmp[1108]*kernel[4]+tmp[1109]*kernel[5]+tmp[1207]*kernel[6]+tmp[1208]*kernel[7]+tmp[1209]*kernel[8];
				ans[1109]<=tmp[1008]*kernel[0]+tmp[1009]*kernel[1]+tmp[1010]*kernel[2]+tmp[1108]*kernel[3]+tmp[1109]*kernel[4]+tmp[1110]*kernel[5]+tmp[1208]*kernel[6]+tmp[1209]*kernel[7]+tmp[1210]*kernel[8];
				ans[1110]<=tmp[1009]*kernel[0]+tmp[1010]*kernel[1]+tmp[1011]*kernel[2]+tmp[1109]*kernel[3]+tmp[1110]*kernel[4]+tmp[1111]*kernel[5]+tmp[1209]*kernel[6]+tmp[1210]*kernel[7]+tmp[1211]*kernel[8];
				ans[1111]<=tmp[1010]*kernel[0]+tmp[1011]*kernel[1]+tmp[1012]*kernel[2]+tmp[1110]*kernel[3]+tmp[1111]*kernel[4]+tmp[1112]*kernel[5]+tmp[1210]*kernel[6]+tmp[1211]*kernel[7]+tmp[1212]*kernel[8];
				ans[1112]<=tmp[1011]*kernel[0]+tmp[1012]*kernel[1]+tmp[1013]*kernel[2]+tmp[1111]*kernel[3]+tmp[1112]*kernel[4]+tmp[1113]*kernel[5]+tmp[1211]*kernel[6]+tmp[1212]*kernel[7]+tmp[1213]*kernel[8];
				ans[1113]<=tmp[1012]*kernel[0]+tmp[1013]*kernel[1]+tmp[1014]*kernel[2]+tmp[1112]*kernel[3]+tmp[1113]*kernel[4]+tmp[1114]*kernel[5]+tmp[1212]*kernel[6]+tmp[1213]*kernel[7]+tmp[1214]*kernel[8];
				ans[1114]<=tmp[1013]*kernel[0]+tmp[1014]*kernel[1]+tmp[1015]*kernel[2]+tmp[1113]*kernel[3]+tmp[1114]*kernel[4]+tmp[1115]*kernel[5]+tmp[1213]*kernel[6]+tmp[1214]*kernel[7]+tmp[1215]*kernel[8];
				ans[1115]<=tmp[1014]*kernel[0]+tmp[1015]*kernel[1]+tmp[1016]*kernel[2]+tmp[1114]*kernel[3]+tmp[1115]*kernel[4]+tmp[1116]*kernel[5]+tmp[1214]*kernel[6]+tmp[1215]*kernel[7]+tmp[1216]*kernel[8];
				ans[1116]<=tmp[1015]*kernel[0]+tmp[1016]*kernel[1]+tmp[1017]*kernel[2]+tmp[1115]*kernel[3]+tmp[1116]*kernel[4]+tmp[1117]*kernel[5]+tmp[1215]*kernel[6]+tmp[1216]*kernel[7]+tmp[1217]*kernel[8];
				ans[1117]<=tmp[1016]*kernel[0]+tmp[1017]*kernel[1]+tmp[1018]*kernel[2]+tmp[1116]*kernel[3]+tmp[1117]*kernel[4]+tmp[1118]*kernel[5]+tmp[1216]*kernel[6]+tmp[1217]*kernel[7]+tmp[1218]*kernel[8];
				ans[1118]<=tmp[1017]*kernel[0]+tmp[1018]*kernel[1]+tmp[1019]*kernel[2]+tmp[1117]*kernel[3]+tmp[1118]*kernel[4]+tmp[1119]*kernel[5]+tmp[1217]*kernel[6]+tmp[1218]*kernel[7]+tmp[1219]*kernel[8];
				ans[1119]<=tmp[1018]*kernel[0]+tmp[1019]*kernel[1]+tmp[1020]*kernel[2]+tmp[1118]*kernel[3]+tmp[1119]*kernel[4]+tmp[1120]*kernel[5]+tmp[1218]*kernel[6]+tmp[1219]*kernel[7]+tmp[1220]*kernel[8];
				ans[1120]<=tmp[1019]*kernel[0]+tmp[1020]*kernel[1]+tmp[1021]*kernel[2]+tmp[1119]*kernel[3]+tmp[1120]*kernel[4]+tmp[1121]*kernel[5]+tmp[1219]*kernel[6]+tmp[1220]*kernel[7]+tmp[1221]*kernel[8];
				ans[1121]<=tmp[1020]*kernel[0]+tmp[1021]*kernel[1]+tmp[1022]*kernel[2]+tmp[1120]*kernel[3]+tmp[1121]*kernel[4]+tmp[1122]*kernel[5]+tmp[1220]*kernel[6]+tmp[1221]*kernel[7]+tmp[1222]*kernel[8];
				ans[1122]<=tmp[1021]*kernel[0]+tmp[1022]*kernel[1]+tmp[1023]*kernel[2]+tmp[1121]*kernel[3]+tmp[1122]*kernel[4]+tmp[1123]*kernel[5]+tmp[1221]*kernel[6]+tmp[1222]*kernel[7]+tmp[1223]*kernel[8];
				ans[1123]<=tmp[1022]*kernel[0]+tmp[1023]*kernel[1]+tmp[1024]*kernel[2]+tmp[1122]*kernel[3]+tmp[1123]*kernel[4]+tmp[1124]*kernel[5]+tmp[1222]*kernel[6]+tmp[1223]*kernel[7]+tmp[1224]*kernel[8];
				ans[1124]<=tmp[1023]*kernel[0]+tmp[1024]*kernel[1]+tmp[1025]*kernel[2]+tmp[1123]*kernel[3]+tmp[1124]*kernel[4]+tmp[1125]*kernel[5]+tmp[1223]*kernel[6]+tmp[1224]*kernel[7]+tmp[1225]*kernel[8];
				ans[1125]<=tmp[1024]*kernel[0]+tmp[1025]*kernel[1]+tmp[1026]*kernel[2]+tmp[1124]*kernel[3]+tmp[1125]*kernel[4]+tmp[1126]*kernel[5]+tmp[1224]*kernel[6]+tmp[1225]*kernel[7]+tmp[1226]*kernel[8];
				ans[1126]<=tmp[1025]*kernel[0]+tmp[1026]*kernel[1]+tmp[1027]*kernel[2]+tmp[1125]*kernel[3]+tmp[1126]*kernel[4]+tmp[1127]*kernel[5]+tmp[1225]*kernel[6]+tmp[1226]*kernel[7]+tmp[1227]*kernel[8];
				ans[1127]<=tmp[1026]*kernel[0]+tmp[1027]*kernel[1]+tmp[1028]*kernel[2]+tmp[1126]*kernel[3]+tmp[1127]*kernel[4]+tmp[1128]*kernel[5]+tmp[1226]*kernel[6]+tmp[1227]*kernel[7]+tmp[1228]*kernel[8];
				ans[1128]<=tmp[1027]*kernel[0]+tmp[1028]*kernel[1]+tmp[1029]*kernel[2]+tmp[1127]*kernel[3]+tmp[1128]*kernel[4]+tmp[1129]*kernel[5]+tmp[1227]*kernel[6]+tmp[1228]*kernel[7]+tmp[1229]*kernel[8];
				ans[1129]<=tmp[1028]*kernel[0]+tmp[1029]*kernel[1]+tmp[1030]*kernel[2]+tmp[1128]*kernel[3]+tmp[1129]*kernel[4]+tmp[1130]*kernel[5]+tmp[1228]*kernel[6]+tmp[1229]*kernel[7]+tmp[1230]*kernel[8];
				ans[1130]<=tmp[1029]*kernel[0]+tmp[1030]*kernel[1]+tmp[1031]*kernel[2]+tmp[1129]*kernel[3]+tmp[1130]*kernel[4]+tmp[1131]*kernel[5]+tmp[1229]*kernel[6]+tmp[1230]*kernel[7]+tmp[1231]*kernel[8];
				ans[1131]<=tmp[1030]*kernel[0]+tmp[1031]*kernel[1]+tmp[1032]*kernel[2]+tmp[1130]*kernel[3]+tmp[1131]*kernel[4]+tmp[1132]*kernel[5]+tmp[1230]*kernel[6]+tmp[1231]*kernel[7]+tmp[1232]*kernel[8];
				ans[1132]<=tmp[1031]*kernel[0]+tmp[1032]*kernel[1]+tmp[1033]*kernel[2]+tmp[1131]*kernel[3]+tmp[1132]*kernel[4]+tmp[1133]*kernel[5]+tmp[1231]*kernel[6]+tmp[1232]*kernel[7]+tmp[1233]*kernel[8];
				ans[1133]<=tmp[1032]*kernel[0]+tmp[1033]*kernel[1]+tmp[1034]*kernel[2]+tmp[1132]*kernel[3]+tmp[1133]*kernel[4]+tmp[1134]*kernel[5]+tmp[1232]*kernel[6]+tmp[1233]*kernel[7]+tmp[1234]*kernel[8];
				ans[1134]<=tmp[1033]*kernel[0]+tmp[1034]*kernel[1]+tmp[1035]*kernel[2]+tmp[1133]*kernel[3]+tmp[1134]*kernel[4]+tmp[1135]*kernel[5]+tmp[1233]*kernel[6]+tmp[1234]*kernel[7]+tmp[1235]*kernel[8];
				ans[1135]<=tmp[1034]*kernel[0]+tmp[1035]*kernel[1]+tmp[1036]*kernel[2]+tmp[1134]*kernel[3]+tmp[1135]*kernel[4]+tmp[1136]*kernel[5]+tmp[1234]*kernel[6]+tmp[1235]*kernel[7]+tmp[1236]*kernel[8];
				ans[1136]<=tmp[1035]*kernel[0]+tmp[1036]*kernel[1]+tmp[1037]*kernel[2]+tmp[1135]*kernel[3]+tmp[1136]*kernel[4]+tmp[1137]*kernel[5]+tmp[1235]*kernel[6]+tmp[1236]*kernel[7]+tmp[1237]*kernel[8];
				ans[1137]<=tmp[1036]*kernel[0]+tmp[1037]*kernel[1]+tmp[1038]*kernel[2]+tmp[1136]*kernel[3]+tmp[1137]*kernel[4]+tmp[1138]*kernel[5]+tmp[1236]*kernel[6]+tmp[1237]*kernel[7]+tmp[1238]*kernel[8];
				ans[1138]<=tmp[1037]*kernel[0]+tmp[1038]*kernel[1]+tmp[1039]*kernel[2]+tmp[1137]*kernel[3]+tmp[1138]*kernel[4]+tmp[1139]*kernel[5]+tmp[1237]*kernel[6]+tmp[1238]*kernel[7]+tmp[1239]*kernel[8];
				ans[1139]<=tmp[1038]*kernel[0]+tmp[1039]*kernel[1]+tmp[1040]*kernel[2]+tmp[1138]*kernel[3]+tmp[1139]*kernel[4]+tmp[1140]*kernel[5]+tmp[1238]*kernel[6]+tmp[1239]*kernel[7]+tmp[1240]*kernel[8];
				ans[1140]<=tmp[1039]*kernel[0]+tmp[1040]*kernel[1]+tmp[1041]*kernel[2]+tmp[1139]*kernel[3]+tmp[1140]*kernel[4]+tmp[1141]*kernel[5]+tmp[1239]*kernel[6]+tmp[1240]*kernel[7]+tmp[1241]*kernel[8];
				ans[1141]<=tmp[1040]*kernel[0]+tmp[1041]*kernel[1]+tmp[1042]*kernel[2]+tmp[1140]*kernel[3]+tmp[1141]*kernel[4]+tmp[1142]*kernel[5]+tmp[1240]*kernel[6]+tmp[1241]*kernel[7]+tmp[1242]*kernel[8];
				ans[1142]<=tmp[1041]*kernel[0]+tmp[1042]*kernel[1]+tmp[1043]*kernel[2]+tmp[1141]*kernel[3]+tmp[1142]*kernel[4]+tmp[1143]*kernel[5]+tmp[1241]*kernel[6]+tmp[1242]*kernel[7]+tmp[1243]*kernel[8];
				ans[1143]<=tmp[1042]*kernel[0]+tmp[1043]*kernel[1]+tmp[1044]*kernel[2]+tmp[1142]*kernel[3]+tmp[1143]*kernel[4]+tmp[1144]*kernel[5]+tmp[1242]*kernel[6]+tmp[1243]*kernel[7]+tmp[1244]*kernel[8];
				ans[1144]<=tmp[1043]*kernel[0]+tmp[1044]*kernel[1]+tmp[1045]*kernel[2]+tmp[1143]*kernel[3]+tmp[1144]*kernel[4]+tmp[1145]*kernel[5]+tmp[1243]*kernel[6]+tmp[1244]*kernel[7]+tmp[1245]*kernel[8];
				ans[1145]<=tmp[1044]*kernel[0]+tmp[1045]*kernel[1]+tmp[1046]*kernel[2]+tmp[1144]*kernel[3]+tmp[1145]*kernel[4]+tmp[1146]*kernel[5]+tmp[1244]*kernel[6]+tmp[1245]*kernel[7]+tmp[1246]*kernel[8];
				ans[1146]<=tmp[1045]*kernel[0]+tmp[1046]*kernel[1]+tmp[1047]*kernel[2]+tmp[1145]*kernel[3]+tmp[1146]*kernel[4]+tmp[1147]*kernel[5]+tmp[1245]*kernel[6]+tmp[1246]*kernel[7]+tmp[1247]*kernel[8];
				ans[1147]<=tmp[1046]*kernel[0]+tmp[1047]*kernel[1]+tmp[1048]*kernel[2]+tmp[1146]*kernel[3]+tmp[1147]*kernel[4]+tmp[1148]*kernel[5]+tmp[1246]*kernel[6]+tmp[1247]*kernel[7]+tmp[1248]*kernel[8];
				ans[1148]<=tmp[1047]*kernel[0]+tmp[1048]*kernel[1]+tmp[1049]*kernel[2]+tmp[1147]*kernel[3]+tmp[1148]*kernel[4]+tmp[1149]*kernel[5]+tmp[1247]*kernel[6]+tmp[1248]*kernel[7]+tmp[1249]*kernel[8];
				ans[1149]<=tmp[1048]*kernel[0]+tmp[1049]*kernel[1]+tmp[1050]*kernel[2]+tmp[1148]*kernel[3]+tmp[1149]*kernel[4]+tmp[1150]*kernel[5]+tmp[1248]*kernel[6]+tmp[1249]*kernel[7]+tmp[1250]*kernel[8];
				ans[1150]<=tmp[1049]*kernel[0]+tmp[1050]*kernel[1]+tmp[1051]*kernel[2]+tmp[1149]*kernel[3]+tmp[1150]*kernel[4]+tmp[1151]*kernel[5]+tmp[1249]*kernel[6]+tmp[1250]*kernel[7]+tmp[1251]*kernel[8];
				ans[1151]<=tmp[1050]*kernel[0]+tmp[1051]*kernel[1]+tmp[1052]*kernel[2]+tmp[1150]*kernel[3]+tmp[1151]*kernel[4]+tmp[1152]*kernel[5]+tmp[1250]*kernel[6]+tmp[1251]*kernel[7]+tmp[1252]*kernel[8];
				ans[1152]<=tmp[1051]*kernel[0]+tmp[1052]*kernel[1]+tmp[1053]*kernel[2]+tmp[1151]*kernel[3]+tmp[1152]*kernel[4]+tmp[1153]*kernel[5]+tmp[1251]*kernel[6]+tmp[1252]*kernel[7]+tmp[1253]*kernel[8];
				ans[1153]<=tmp[1052]*kernel[0]+tmp[1053]*kernel[1]+tmp[1054]*kernel[2]+tmp[1152]*kernel[3]+tmp[1153]*kernel[4]+tmp[1154]*kernel[5]+tmp[1252]*kernel[6]+tmp[1253]*kernel[7]+tmp[1254]*kernel[8];
				ans[1154]<=tmp[1053]*kernel[0]+tmp[1054]*kernel[1]+tmp[1055]*kernel[2]+tmp[1153]*kernel[3]+tmp[1154]*kernel[4]+tmp[1155]*kernel[5]+tmp[1253]*kernel[6]+tmp[1254]*kernel[7]+tmp[1255]*kernel[8];
				ans[1155]<=tmp[1054]*kernel[0]+tmp[1055]*kernel[1]+tmp[1056]*kernel[2]+tmp[1154]*kernel[3]+tmp[1155]*kernel[4]+tmp[1156]*kernel[5]+tmp[1254]*kernel[6]+tmp[1255]*kernel[7]+tmp[1256]*kernel[8];
				ans[1156]<=tmp[1055]*kernel[0]+tmp[1056]*kernel[1]+tmp[1057]*kernel[2]+tmp[1155]*kernel[3]+tmp[1156]*kernel[4]+tmp[1157]*kernel[5]+tmp[1255]*kernel[6]+tmp[1256]*kernel[7]+tmp[1257]*kernel[8];
				ans[1157]<=tmp[1056]*kernel[0]+tmp[1057]*kernel[1]+tmp[1058]*kernel[2]+tmp[1156]*kernel[3]+tmp[1157]*kernel[4]+tmp[1158]*kernel[5]+tmp[1256]*kernel[6]+tmp[1257]*kernel[7]+tmp[1258]*kernel[8];
				ans[1158]<=tmp[1057]*kernel[0]+tmp[1058]*kernel[1]+tmp[1059]*kernel[2]+tmp[1157]*kernel[3]+tmp[1158]*kernel[4]+tmp[1159]*kernel[5]+tmp[1257]*kernel[6]+tmp[1258]*kernel[7]+tmp[1259]*kernel[8];
				ans[1159]<=tmp[1058]*kernel[0]+tmp[1059]*kernel[1]+tmp[1060]*kernel[2]+tmp[1158]*kernel[3]+tmp[1159]*kernel[4]+tmp[1160]*kernel[5]+tmp[1258]*kernel[6]+tmp[1259]*kernel[7]+tmp[1260]*kernel[8];
				ans[1160]<=tmp[1059]*kernel[0]+tmp[1060]*kernel[1]+tmp[1061]*kernel[2]+tmp[1159]*kernel[3]+tmp[1160]*kernel[4]+tmp[1161]*kernel[5]+tmp[1259]*kernel[6]+tmp[1260]*kernel[7]+tmp[1261]*kernel[8];
				ans[1161]<=tmp[1060]*kernel[0]+tmp[1061]*kernel[1]+tmp[1062]*kernel[2]+tmp[1160]*kernel[3]+tmp[1161]*kernel[4]+tmp[1162]*kernel[5]+tmp[1260]*kernel[6]+tmp[1261]*kernel[7]+tmp[1262]*kernel[8];
				ans[1162]<=tmp[1061]*kernel[0]+tmp[1062]*kernel[1]+tmp[1063]*kernel[2]+tmp[1161]*kernel[3]+tmp[1162]*kernel[4]+tmp[1163]*kernel[5]+tmp[1261]*kernel[6]+tmp[1262]*kernel[7]+tmp[1263]*kernel[8];
				ans[1163]<=tmp[1062]*kernel[0]+tmp[1063]*kernel[1]+tmp[1064]*kernel[2]+tmp[1162]*kernel[3]+tmp[1163]*kernel[4]+tmp[1164]*kernel[5]+tmp[1262]*kernel[6]+tmp[1263]*kernel[7]+tmp[1264]*kernel[8];
				ans[1164]<=tmp[1063]*kernel[0]+tmp[1064]*kernel[1]+tmp[1065]*kernel[2]+tmp[1163]*kernel[3]+tmp[1164]*kernel[4]+tmp[1165]*kernel[5]+tmp[1263]*kernel[6]+tmp[1264]*kernel[7]+tmp[1265]*kernel[8];
				ans[1165]<=tmp[1064]*kernel[0]+tmp[1065]*kernel[1]+tmp[1066]*kernel[2]+tmp[1164]*kernel[3]+tmp[1165]*kernel[4]+tmp[1166]*kernel[5]+tmp[1264]*kernel[6]+tmp[1265]*kernel[7]+tmp[1266]*kernel[8];
				ans[1166]<=tmp[1065]*kernel[0]+tmp[1066]*kernel[1]+tmp[1067]*kernel[2]+tmp[1165]*kernel[3]+tmp[1166]*kernel[4]+tmp[1167]*kernel[5]+tmp[1265]*kernel[6]+tmp[1266]*kernel[7]+tmp[1267]*kernel[8];
				ans[1167]<=tmp[1066]*kernel[0]+tmp[1067]*kernel[1]+tmp[1068]*kernel[2]+tmp[1166]*kernel[3]+tmp[1167]*kernel[4]+tmp[1168]*kernel[5]+tmp[1266]*kernel[6]+tmp[1267]*kernel[7]+tmp[1268]*kernel[8];
				ans[1168]<=tmp[1067]*kernel[0]+tmp[1068]*kernel[1]+tmp[1069]*kernel[2]+tmp[1167]*kernel[3]+tmp[1168]*kernel[4]+tmp[1169]*kernel[5]+tmp[1267]*kernel[6]+tmp[1268]*kernel[7]+tmp[1269]*kernel[8];
				ans[1169]<=tmp[1068]*kernel[0]+tmp[1069]*kernel[1]+tmp[1070]*kernel[2]+tmp[1168]*kernel[3]+tmp[1169]*kernel[4]+tmp[1170]*kernel[5]+tmp[1268]*kernel[6]+tmp[1269]*kernel[7]+tmp[1270]*kernel[8];
				ans[1170]<=tmp[1069]*kernel[0]+tmp[1070]*kernel[1]+tmp[1071]*kernel[2]+tmp[1169]*kernel[3]+tmp[1170]*kernel[4]+tmp[1171]*kernel[5]+tmp[1269]*kernel[6]+tmp[1270]*kernel[7]+tmp[1271]*kernel[8];
				ans[1171]<=tmp[1070]*kernel[0]+tmp[1071]*kernel[1]+tmp[1072]*kernel[2]+tmp[1170]*kernel[3]+tmp[1171]*kernel[4]+tmp[1172]*kernel[5]+tmp[1270]*kernel[6]+tmp[1271]*kernel[7]+tmp[1272]*kernel[8];
				ans[1172]<=tmp[1071]*kernel[0]+tmp[1072]*kernel[1]+tmp[1073]*kernel[2]+tmp[1171]*kernel[3]+tmp[1172]*kernel[4]+tmp[1173]*kernel[5]+tmp[1271]*kernel[6]+tmp[1272]*kernel[7]+tmp[1273]*kernel[8];
				ans[1173]<=tmp[1072]*kernel[0]+tmp[1073]*kernel[1]+tmp[1074]*kernel[2]+tmp[1172]*kernel[3]+tmp[1173]*kernel[4]+tmp[1174]*kernel[5]+tmp[1272]*kernel[6]+tmp[1273]*kernel[7]+tmp[1274]*kernel[8];
				ans[1174]<=tmp[1073]*kernel[0]+tmp[1074]*kernel[1]+tmp[1075]*kernel[2]+tmp[1173]*kernel[3]+tmp[1174]*kernel[4]+tmp[1175]*kernel[5]+tmp[1273]*kernel[6]+tmp[1274]*kernel[7]+tmp[1275]*kernel[8];
				ans[1175]<=tmp[1074]*kernel[0]+tmp[1075]*kernel[1]+tmp[1076]*kernel[2]+tmp[1174]*kernel[3]+tmp[1175]*kernel[4]+tmp[1176]*kernel[5]+tmp[1274]*kernel[6]+tmp[1275]*kernel[7]+tmp[1276]*kernel[8];
				ans[1176]<=tmp[1075]*kernel[0]+tmp[1076]*kernel[1]+tmp[1077]*kernel[2]+tmp[1175]*kernel[3]+tmp[1176]*kernel[4]+tmp[1177]*kernel[5]+tmp[1275]*kernel[6]+tmp[1276]*kernel[7]+tmp[1277]*kernel[8];
				ans[1177]<=tmp[1076]*kernel[0]+tmp[1077]*kernel[1]+tmp[1078]*kernel[2]+tmp[1176]*kernel[3]+tmp[1177]*kernel[4]+tmp[1178]*kernel[5]+tmp[1276]*kernel[6]+tmp[1277]*kernel[7]+tmp[1278]*kernel[8];
				ans[1178]<=tmp[1077]*kernel[0]+tmp[1078]*kernel[1]+tmp[1079]*kernel[2]+tmp[1177]*kernel[3]+tmp[1178]*kernel[4]+tmp[1179]*kernel[5]+tmp[1277]*kernel[6]+tmp[1278]*kernel[7]+tmp[1279]*kernel[8];
				ans[1179]<=tmp[1078]*kernel[0]+tmp[1079]*kernel[1]+tmp[1080]*kernel[2]+tmp[1178]*kernel[3]+tmp[1179]*kernel[4]+tmp[1180]*kernel[5]+tmp[1278]*kernel[6]+tmp[1279]*kernel[7]+tmp[1280]*kernel[8];
				ans[1180]<=tmp[1079]*kernel[0]+tmp[1080]*kernel[1]+tmp[1081]*kernel[2]+tmp[1179]*kernel[3]+tmp[1180]*kernel[4]+tmp[1181]*kernel[5]+tmp[1279]*kernel[6]+tmp[1280]*kernel[7]+tmp[1281]*kernel[8];
				ans[1181]<=tmp[1080]*kernel[0]+tmp[1081]*kernel[1]+tmp[1082]*kernel[2]+tmp[1180]*kernel[3]+tmp[1181]*kernel[4]+tmp[1182]*kernel[5]+tmp[1280]*kernel[6]+tmp[1281]*kernel[7]+tmp[1282]*kernel[8];
				ans[1182]<=tmp[1081]*kernel[0]+tmp[1082]*kernel[1]+tmp[1083]*kernel[2]+tmp[1181]*kernel[3]+tmp[1182]*kernel[4]+tmp[1183]*kernel[5]+tmp[1281]*kernel[6]+tmp[1282]*kernel[7]+tmp[1283]*kernel[8];
				ans[1183]<=tmp[1082]*kernel[0]+tmp[1083]*kernel[1]+tmp[1084]*kernel[2]+tmp[1182]*kernel[3]+tmp[1183]*kernel[4]+tmp[1184]*kernel[5]+tmp[1282]*kernel[6]+tmp[1283]*kernel[7]+tmp[1284]*kernel[8];
				ans[1184]<=tmp[1083]*kernel[0]+tmp[1084]*kernel[1]+tmp[1085]*kernel[2]+tmp[1183]*kernel[3]+tmp[1184]*kernel[4]+tmp[1185]*kernel[5]+tmp[1283]*kernel[6]+tmp[1284]*kernel[7]+tmp[1285]*kernel[8];
				ans[1185]<=tmp[1084]*kernel[0]+tmp[1085]*kernel[1]+tmp[1086]*kernel[2]+tmp[1184]*kernel[3]+tmp[1185]*kernel[4]+tmp[1186]*kernel[5]+tmp[1284]*kernel[6]+tmp[1285]*kernel[7]+tmp[1286]*kernel[8];
				ans[1186]<=tmp[1085]*kernel[0]+tmp[1086]*kernel[1]+tmp[1087]*kernel[2]+tmp[1185]*kernel[3]+tmp[1186]*kernel[4]+tmp[1187]*kernel[5]+tmp[1285]*kernel[6]+tmp[1286]*kernel[7]+tmp[1287]*kernel[8];
				ans[1187]<=tmp[1086]*kernel[0]+tmp[1087]*kernel[1]+tmp[1088]*kernel[2]+tmp[1186]*kernel[3]+tmp[1187]*kernel[4]+tmp[1188]*kernel[5]+tmp[1286]*kernel[6]+tmp[1287]*kernel[7]+tmp[1288]*kernel[8];
				ans[1188]<=tmp[1087]*kernel[0]+tmp[1088]*kernel[1]+tmp[1089]*kernel[2]+tmp[1187]*kernel[3]+tmp[1188]*kernel[4]+tmp[1189]*kernel[5]+tmp[1287]*kernel[6]+tmp[1288]*kernel[7]+tmp[1289]*kernel[8];
				ans[1189]<=tmp[1088]*kernel[0]+tmp[1089]*kernel[1]+tmp[1090]*kernel[2]+tmp[1188]*kernel[3]+tmp[1189]*kernel[4]+tmp[1190]*kernel[5]+tmp[1288]*kernel[6]+tmp[1289]*kernel[7]+tmp[1290]*kernel[8];
				ans[1190]<=tmp[1089]*kernel[0]+tmp[1090]*kernel[1]+tmp[1091]*kernel[2]+tmp[1189]*kernel[3]+tmp[1190]*kernel[4]+tmp[1191]*kernel[5]+tmp[1289]*kernel[6]+tmp[1290]*kernel[7]+tmp[1291]*kernel[8];
				ans[1191]<=tmp[1090]*kernel[0]+tmp[1091]*kernel[1]+tmp[1092]*kernel[2]+tmp[1190]*kernel[3]+tmp[1191]*kernel[4]+tmp[1192]*kernel[5]+tmp[1290]*kernel[6]+tmp[1291]*kernel[7]+tmp[1292]*kernel[8];
				ans[1192]<=tmp[1091]*kernel[0]+tmp[1092]*kernel[1]+tmp[1093]*kernel[2]+tmp[1191]*kernel[3]+tmp[1192]*kernel[4]+tmp[1193]*kernel[5]+tmp[1291]*kernel[6]+tmp[1292]*kernel[7]+tmp[1293]*kernel[8];
				ans[1193]<=tmp[1092]*kernel[0]+tmp[1093]*kernel[1]+tmp[1094]*kernel[2]+tmp[1192]*kernel[3]+tmp[1193]*kernel[4]+tmp[1194]*kernel[5]+tmp[1292]*kernel[6]+tmp[1293]*kernel[7]+tmp[1294]*kernel[8];
				ans[1194]<=tmp[1093]*kernel[0]+tmp[1094]*kernel[1]+tmp[1095]*kernel[2]+tmp[1193]*kernel[3]+tmp[1194]*kernel[4]+tmp[1195]*kernel[5]+tmp[1293]*kernel[6]+tmp[1294]*kernel[7]+tmp[1295]*kernel[8];
				ans[1195]<=tmp[1094]*kernel[0]+tmp[1095]*kernel[1]+tmp[1096]*kernel[2]+tmp[1194]*kernel[3]+tmp[1195]*kernel[4]+tmp[1196]*kernel[5]+tmp[1294]*kernel[6]+tmp[1295]*kernel[7]+tmp[1296]*kernel[8];
				ans[1196]<=tmp[1095]*kernel[0]+tmp[1096]*kernel[1]+tmp[1097]*kernel[2]+tmp[1195]*kernel[3]+tmp[1196]*kernel[4]+tmp[1197]*kernel[5]+tmp[1295]*kernel[6]+tmp[1296]*kernel[7]+tmp[1297]*kernel[8];
				ans[1197]<=tmp[1096]*kernel[0]+tmp[1097]*kernel[1]+tmp[1098]*kernel[2]+tmp[1196]*kernel[3]+tmp[1197]*kernel[4]+tmp[1198]*kernel[5]+tmp[1296]*kernel[6]+tmp[1297]*kernel[7]+tmp[1298]*kernel[8];
				ans[1198]<=tmp[1097]*kernel[0]+tmp[1098]*kernel[1]+tmp[1099]*kernel[2]+tmp[1197]*kernel[3]+tmp[1198]*kernel[4]+tmp[1199]*kernel[5]+tmp[1297]*kernel[6]+tmp[1298]*kernel[7]+tmp[1299]*kernel[8];
				ans[1199]<=tmp[1098]*kernel[0]+tmp[1099]*kernel[1]+tmp[1198]*kernel[3]+tmp[1199]*kernel[4]+tmp[1298]*kernel[6]+tmp[1299]*kernel[7];
				ans[1200]<=tmp[1100]*kernel[1]+tmp[1101]*kernel[2]+tmp[1200]*kernel[4]+tmp[1201]*kernel[5]+tmp[1300]*kernel[7]+tmp[1301]*kernel[8];
				ans[1201]<=tmp[1100]*kernel[0]+tmp[1101]*kernel[1]+tmp[1102]*kernel[2]+tmp[1200]*kernel[3]+tmp[1201]*kernel[4]+tmp[1202]*kernel[5]+tmp[1300]*kernel[6]+tmp[1301]*kernel[7]+tmp[1302]*kernel[8];
				ans[1202]<=tmp[1101]*kernel[0]+tmp[1102]*kernel[1]+tmp[1103]*kernel[2]+tmp[1201]*kernel[3]+tmp[1202]*kernel[4]+tmp[1203]*kernel[5]+tmp[1301]*kernel[6]+tmp[1302]*kernel[7]+tmp[1303]*kernel[8];
				ans[1203]<=tmp[1102]*kernel[0]+tmp[1103]*kernel[1]+tmp[1104]*kernel[2]+tmp[1202]*kernel[3]+tmp[1203]*kernel[4]+tmp[1204]*kernel[5]+tmp[1302]*kernel[6]+tmp[1303]*kernel[7]+tmp[1304]*kernel[8];
				ans[1204]<=tmp[1103]*kernel[0]+tmp[1104]*kernel[1]+tmp[1105]*kernel[2]+tmp[1203]*kernel[3]+tmp[1204]*kernel[4]+tmp[1205]*kernel[5]+tmp[1303]*kernel[6]+tmp[1304]*kernel[7]+tmp[1305]*kernel[8];
				ans[1205]<=tmp[1104]*kernel[0]+tmp[1105]*kernel[1]+tmp[1106]*kernel[2]+tmp[1204]*kernel[3]+tmp[1205]*kernel[4]+tmp[1206]*kernel[5]+tmp[1304]*kernel[6]+tmp[1305]*kernel[7]+tmp[1306]*kernel[8];
				ans[1206]<=tmp[1105]*kernel[0]+tmp[1106]*kernel[1]+tmp[1107]*kernel[2]+tmp[1205]*kernel[3]+tmp[1206]*kernel[4]+tmp[1207]*kernel[5]+tmp[1305]*kernel[6]+tmp[1306]*kernel[7]+tmp[1307]*kernel[8];
				ans[1207]<=tmp[1106]*kernel[0]+tmp[1107]*kernel[1]+tmp[1108]*kernel[2]+tmp[1206]*kernel[3]+tmp[1207]*kernel[4]+tmp[1208]*kernel[5]+tmp[1306]*kernel[6]+tmp[1307]*kernel[7]+tmp[1308]*kernel[8];
				ans[1208]<=tmp[1107]*kernel[0]+tmp[1108]*kernel[1]+tmp[1109]*kernel[2]+tmp[1207]*kernel[3]+tmp[1208]*kernel[4]+tmp[1209]*kernel[5]+tmp[1307]*kernel[6]+tmp[1308]*kernel[7]+tmp[1309]*kernel[8];
				ans[1209]<=tmp[1108]*kernel[0]+tmp[1109]*kernel[1]+tmp[1110]*kernel[2]+tmp[1208]*kernel[3]+tmp[1209]*kernel[4]+tmp[1210]*kernel[5]+tmp[1308]*kernel[6]+tmp[1309]*kernel[7]+tmp[1310]*kernel[8];
				ans[1210]<=tmp[1109]*kernel[0]+tmp[1110]*kernel[1]+tmp[1111]*kernel[2]+tmp[1209]*kernel[3]+tmp[1210]*kernel[4]+tmp[1211]*kernel[5]+tmp[1309]*kernel[6]+tmp[1310]*kernel[7]+tmp[1311]*kernel[8];
				ans[1211]<=tmp[1110]*kernel[0]+tmp[1111]*kernel[1]+tmp[1112]*kernel[2]+tmp[1210]*kernel[3]+tmp[1211]*kernel[4]+tmp[1212]*kernel[5]+tmp[1310]*kernel[6]+tmp[1311]*kernel[7]+tmp[1312]*kernel[8];
				ans[1212]<=tmp[1111]*kernel[0]+tmp[1112]*kernel[1]+tmp[1113]*kernel[2]+tmp[1211]*kernel[3]+tmp[1212]*kernel[4]+tmp[1213]*kernel[5]+tmp[1311]*kernel[6]+tmp[1312]*kernel[7]+tmp[1313]*kernel[8];
				ans[1213]<=tmp[1112]*kernel[0]+tmp[1113]*kernel[1]+tmp[1114]*kernel[2]+tmp[1212]*kernel[3]+tmp[1213]*kernel[4]+tmp[1214]*kernel[5]+tmp[1312]*kernel[6]+tmp[1313]*kernel[7]+tmp[1314]*kernel[8];
				ans[1214]<=tmp[1113]*kernel[0]+tmp[1114]*kernel[1]+tmp[1115]*kernel[2]+tmp[1213]*kernel[3]+tmp[1214]*kernel[4]+tmp[1215]*kernel[5]+tmp[1313]*kernel[6]+tmp[1314]*kernel[7]+tmp[1315]*kernel[8];
				ans[1215]<=tmp[1114]*kernel[0]+tmp[1115]*kernel[1]+tmp[1116]*kernel[2]+tmp[1214]*kernel[3]+tmp[1215]*kernel[4]+tmp[1216]*kernel[5]+tmp[1314]*kernel[6]+tmp[1315]*kernel[7]+tmp[1316]*kernel[8];
				ans[1216]<=tmp[1115]*kernel[0]+tmp[1116]*kernel[1]+tmp[1117]*kernel[2]+tmp[1215]*kernel[3]+tmp[1216]*kernel[4]+tmp[1217]*kernel[5]+tmp[1315]*kernel[6]+tmp[1316]*kernel[7]+tmp[1317]*kernel[8];
				ans[1217]<=tmp[1116]*kernel[0]+tmp[1117]*kernel[1]+tmp[1118]*kernel[2]+tmp[1216]*kernel[3]+tmp[1217]*kernel[4]+tmp[1218]*kernel[5]+tmp[1316]*kernel[6]+tmp[1317]*kernel[7]+tmp[1318]*kernel[8];
				ans[1218]<=tmp[1117]*kernel[0]+tmp[1118]*kernel[1]+tmp[1119]*kernel[2]+tmp[1217]*kernel[3]+tmp[1218]*kernel[4]+tmp[1219]*kernel[5]+tmp[1317]*kernel[6]+tmp[1318]*kernel[7]+tmp[1319]*kernel[8];
				ans[1219]<=tmp[1118]*kernel[0]+tmp[1119]*kernel[1]+tmp[1120]*kernel[2]+tmp[1218]*kernel[3]+tmp[1219]*kernel[4]+tmp[1220]*kernel[5]+tmp[1318]*kernel[6]+tmp[1319]*kernel[7]+tmp[1320]*kernel[8];
				ans[1220]<=tmp[1119]*kernel[0]+tmp[1120]*kernel[1]+tmp[1121]*kernel[2]+tmp[1219]*kernel[3]+tmp[1220]*kernel[4]+tmp[1221]*kernel[5]+tmp[1319]*kernel[6]+tmp[1320]*kernel[7]+tmp[1321]*kernel[8];
				ans[1221]<=tmp[1120]*kernel[0]+tmp[1121]*kernel[1]+tmp[1122]*kernel[2]+tmp[1220]*kernel[3]+tmp[1221]*kernel[4]+tmp[1222]*kernel[5]+tmp[1320]*kernel[6]+tmp[1321]*kernel[7]+tmp[1322]*kernel[8];
				ans[1222]<=tmp[1121]*kernel[0]+tmp[1122]*kernel[1]+tmp[1123]*kernel[2]+tmp[1221]*kernel[3]+tmp[1222]*kernel[4]+tmp[1223]*kernel[5]+tmp[1321]*kernel[6]+tmp[1322]*kernel[7]+tmp[1323]*kernel[8];
				ans[1223]<=tmp[1122]*kernel[0]+tmp[1123]*kernel[1]+tmp[1124]*kernel[2]+tmp[1222]*kernel[3]+tmp[1223]*kernel[4]+tmp[1224]*kernel[5]+tmp[1322]*kernel[6]+tmp[1323]*kernel[7]+tmp[1324]*kernel[8];
				ans[1224]<=tmp[1123]*kernel[0]+tmp[1124]*kernel[1]+tmp[1125]*kernel[2]+tmp[1223]*kernel[3]+tmp[1224]*kernel[4]+tmp[1225]*kernel[5]+tmp[1323]*kernel[6]+tmp[1324]*kernel[7]+tmp[1325]*kernel[8];
				ans[1225]<=tmp[1124]*kernel[0]+tmp[1125]*kernel[1]+tmp[1126]*kernel[2]+tmp[1224]*kernel[3]+tmp[1225]*kernel[4]+tmp[1226]*kernel[5]+tmp[1324]*kernel[6]+tmp[1325]*kernel[7]+tmp[1326]*kernel[8];
				ans[1226]<=tmp[1125]*kernel[0]+tmp[1126]*kernel[1]+tmp[1127]*kernel[2]+tmp[1225]*kernel[3]+tmp[1226]*kernel[4]+tmp[1227]*kernel[5]+tmp[1325]*kernel[6]+tmp[1326]*kernel[7]+tmp[1327]*kernel[8];
				ans[1227]<=tmp[1126]*kernel[0]+tmp[1127]*kernel[1]+tmp[1128]*kernel[2]+tmp[1226]*kernel[3]+tmp[1227]*kernel[4]+tmp[1228]*kernel[5]+tmp[1326]*kernel[6]+tmp[1327]*kernel[7]+tmp[1328]*kernel[8];
				ans[1228]<=tmp[1127]*kernel[0]+tmp[1128]*kernel[1]+tmp[1129]*kernel[2]+tmp[1227]*kernel[3]+tmp[1228]*kernel[4]+tmp[1229]*kernel[5]+tmp[1327]*kernel[6]+tmp[1328]*kernel[7]+tmp[1329]*kernel[8];
				ans[1229]<=tmp[1128]*kernel[0]+tmp[1129]*kernel[1]+tmp[1130]*kernel[2]+tmp[1228]*kernel[3]+tmp[1229]*kernel[4]+tmp[1230]*kernel[5]+tmp[1328]*kernel[6]+tmp[1329]*kernel[7]+tmp[1330]*kernel[8];
				ans[1230]<=tmp[1129]*kernel[0]+tmp[1130]*kernel[1]+tmp[1131]*kernel[2]+tmp[1229]*kernel[3]+tmp[1230]*kernel[4]+tmp[1231]*kernel[5]+tmp[1329]*kernel[6]+tmp[1330]*kernel[7]+tmp[1331]*kernel[8];
				ans[1231]<=tmp[1130]*kernel[0]+tmp[1131]*kernel[1]+tmp[1132]*kernel[2]+tmp[1230]*kernel[3]+tmp[1231]*kernel[4]+tmp[1232]*kernel[5]+tmp[1330]*kernel[6]+tmp[1331]*kernel[7]+tmp[1332]*kernel[8];
				ans[1232]<=tmp[1131]*kernel[0]+tmp[1132]*kernel[1]+tmp[1133]*kernel[2]+tmp[1231]*kernel[3]+tmp[1232]*kernel[4]+tmp[1233]*kernel[5]+tmp[1331]*kernel[6]+tmp[1332]*kernel[7]+tmp[1333]*kernel[8];
				ans[1233]<=tmp[1132]*kernel[0]+tmp[1133]*kernel[1]+tmp[1134]*kernel[2]+tmp[1232]*kernel[3]+tmp[1233]*kernel[4]+tmp[1234]*kernel[5]+tmp[1332]*kernel[6]+tmp[1333]*kernel[7]+tmp[1334]*kernel[8];
				ans[1234]<=tmp[1133]*kernel[0]+tmp[1134]*kernel[1]+tmp[1135]*kernel[2]+tmp[1233]*kernel[3]+tmp[1234]*kernel[4]+tmp[1235]*kernel[5]+tmp[1333]*kernel[6]+tmp[1334]*kernel[7]+tmp[1335]*kernel[8];
				ans[1235]<=tmp[1134]*kernel[0]+tmp[1135]*kernel[1]+tmp[1136]*kernel[2]+tmp[1234]*kernel[3]+tmp[1235]*kernel[4]+tmp[1236]*kernel[5]+tmp[1334]*kernel[6]+tmp[1335]*kernel[7]+tmp[1336]*kernel[8];
				ans[1236]<=tmp[1135]*kernel[0]+tmp[1136]*kernel[1]+tmp[1137]*kernel[2]+tmp[1235]*kernel[3]+tmp[1236]*kernel[4]+tmp[1237]*kernel[5]+tmp[1335]*kernel[6]+tmp[1336]*kernel[7]+tmp[1337]*kernel[8];
				ans[1237]<=tmp[1136]*kernel[0]+tmp[1137]*kernel[1]+tmp[1138]*kernel[2]+tmp[1236]*kernel[3]+tmp[1237]*kernel[4]+tmp[1238]*kernel[5]+tmp[1336]*kernel[6]+tmp[1337]*kernel[7]+tmp[1338]*kernel[8];
				ans[1238]<=tmp[1137]*kernel[0]+tmp[1138]*kernel[1]+tmp[1139]*kernel[2]+tmp[1237]*kernel[3]+tmp[1238]*kernel[4]+tmp[1239]*kernel[5]+tmp[1337]*kernel[6]+tmp[1338]*kernel[7]+tmp[1339]*kernel[8];
				ans[1239]<=tmp[1138]*kernel[0]+tmp[1139]*kernel[1]+tmp[1140]*kernel[2]+tmp[1238]*kernel[3]+tmp[1239]*kernel[4]+tmp[1240]*kernel[5]+tmp[1338]*kernel[6]+tmp[1339]*kernel[7]+tmp[1340]*kernel[8];
				ans[1240]<=tmp[1139]*kernel[0]+tmp[1140]*kernel[1]+tmp[1141]*kernel[2]+tmp[1239]*kernel[3]+tmp[1240]*kernel[4]+tmp[1241]*kernel[5]+tmp[1339]*kernel[6]+tmp[1340]*kernel[7]+tmp[1341]*kernel[8];
				ans[1241]<=tmp[1140]*kernel[0]+tmp[1141]*kernel[1]+tmp[1142]*kernel[2]+tmp[1240]*kernel[3]+tmp[1241]*kernel[4]+tmp[1242]*kernel[5]+tmp[1340]*kernel[6]+tmp[1341]*kernel[7]+tmp[1342]*kernel[8];
				ans[1242]<=tmp[1141]*kernel[0]+tmp[1142]*kernel[1]+tmp[1143]*kernel[2]+tmp[1241]*kernel[3]+tmp[1242]*kernel[4]+tmp[1243]*kernel[5]+tmp[1341]*kernel[6]+tmp[1342]*kernel[7]+tmp[1343]*kernel[8];
				ans[1243]<=tmp[1142]*kernel[0]+tmp[1143]*kernel[1]+tmp[1144]*kernel[2]+tmp[1242]*kernel[3]+tmp[1243]*kernel[4]+tmp[1244]*kernel[5]+tmp[1342]*kernel[6]+tmp[1343]*kernel[7]+tmp[1344]*kernel[8];
				ans[1244]<=tmp[1143]*kernel[0]+tmp[1144]*kernel[1]+tmp[1145]*kernel[2]+tmp[1243]*kernel[3]+tmp[1244]*kernel[4]+tmp[1245]*kernel[5]+tmp[1343]*kernel[6]+tmp[1344]*kernel[7]+tmp[1345]*kernel[8];
				ans[1245]<=tmp[1144]*kernel[0]+tmp[1145]*kernel[1]+tmp[1146]*kernel[2]+tmp[1244]*kernel[3]+tmp[1245]*kernel[4]+tmp[1246]*kernel[5]+tmp[1344]*kernel[6]+tmp[1345]*kernel[7]+tmp[1346]*kernel[8];
				ans[1246]<=tmp[1145]*kernel[0]+tmp[1146]*kernel[1]+tmp[1147]*kernel[2]+tmp[1245]*kernel[3]+tmp[1246]*kernel[4]+tmp[1247]*kernel[5]+tmp[1345]*kernel[6]+tmp[1346]*kernel[7]+tmp[1347]*kernel[8];
				ans[1247]<=tmp[1146]*kernel[0]+tmp[1147]*kernel[1]+tmp[1148]*kernel[2]+tmp[1246]*kernel[3]+tmp[1247]*kernel[4]+tmp[1248]*kernel[5]+tmp[1346]*kernel[6]+tmp[1347]*kernel[7]+tmp[1348]*kernel[8];
				ans[1248]<=tmp[1147]*kernel[0]+tmp[1148]*kernel[1]+tmp[1149]*kernel[2]+tmp[1247]*kernel[3]+tmp[1248]*kernel[4]+tmp[1249]*kernel[5]+tmp[1347]*kernel[6]+tmp[1348]*kernel[7]+tmp[1349]*kernel[8];
				ans[1249]<=tmp[1148]*kernel[0]+tmp[1149]*kernel[1]+tmp[1150]*kernel[2]+tmp[1248]*kernel[3]+tmp[1249]*kernel[4]+tmp[1250]*kernel[5]+tmp[1348]*kernel[6]+tmp[1349]*kernel[7]+tmp[1350]*kernel[8];
				ans[1250]<=tmp[1149]*kernel[0]+tmp[1150]*kernel[1]+tmp[1151]*kernel[2]+tmp[1249]*kernel[3]+tmp[1250]*kernel[4]+tmp[1251]*kernel[5]+tmp[1349]*kernel[6]+tmp[1350]*kernel[7]+tmp[1351]*kernel[8];
				ans[1251]<=tmp[1150]*kernel[0]+tmp[1151]*kernel[1]+tmp[1152]*kernel[2]+tmp[1250]*kernel[3]+tmp[1251]*kernel[4]+tmp[1252]*kernel[5]+tmp[1350]*kernel[6]+tmp[1351]*kernel[7]+tmp[1352]*kernel[8];
				ans[1252]<=tmp[1151]*kernel[0]+tmp[1152]*kernel[1]+tmp[1153]*kernel[2]+tmp[1251]*kernel[3]+tmp[1252]*kernel[4]+tmp[1253]*kernel[5]+tmp[1351]*kernel[6]+tmp[1352]*kernel[7]+tmp[1353]*kernel[8];
				ans[1253]<=tmp[1152]*kernel[0]+tmp[1153]*kernel[1]+tmp[1154]*kernel[2]+tmp[1252]*kernel[3]+tmp[1253]*kernel[4]+tmp[1254]*kernel[5]+tmp[1352]*kernel[6]+tmp[1353]*kernel[7]+tmp[1354]*kernel[8];
				ans[1254]<=tmp[1153]*kernel[0]+tmp[1154]*kernel[1]+tmp[1155]*kernel[2]+tmp[1253]*kernel[3]+tmp[1254]*kernel[4]+tmp[1255]*kernel[5]+tmp[1353]*kernel[6]+tmp[1354]*kernel[7]+tmp[1355]*kernel[8];
				ans[1255]<=tmp[1154]*kernel[0]+tmp[1155]*kernel[1]+tmp[1156]*kernel[2]+tmp[1254]*kernel[3]+tmp[1255]*kernel[4]+tmp[1256]*kernel[5]+tmp[1354]*kernel[6]+tmp[1355]*kernel[7]+tmp[1356]*kernel[8];
				ans[1256]<=tmp[1155]*kernel[0]+tmp[1156]*kernel[1]+tmp[1157]*kernel[2]+tmp[1255]*kernel[3]+tmp[1256]*kernel[4]+tmp[1257]*kernel[5]+tmp[1355]*kernel[6]+tmp[1356]*kernel[7]+tmp[1357]*kernel[8];
				ans[1257]<=tmp[1156]*kernel[0]+tmp[1157]*kernel[1]+tmp[1158]*kernel[2]+tmp[1256]*kernel[3]+tmp[1257]*kernel[4]+tmp[1258]*kernel[5]+tmp[1356]*kernel[6]+tmp[1357]*kernel[7]+tmp[1358]*kernel[8];
				ans[1258]<=tmp[1157]*kernel[0]+tmp[1158]*kernel[1]+tmp[1159]*kernel[2]+tmp[1257]*kernel[3]+tmp[1258]*kernel[4]+tmp[1259]*kernel[5]+tmp[1357]*kernel[6]+tmp[1358]*kernel[7]+tmp[1359]*kernel[8];
				ans[1259]<=tmp[1158]*kernel[0]+tmp[1159]*kernel[1]+tmp[1160]*kernel[2]+tmp[1258]*kernel[3]+tmp[1259]*kernel[4]+tmp[1260]*kernel[5]+tmp[1358]*kernel[6]+tmp[1359]*kernel[7]+tmp[1360]*kernel[8];
				ans[1260]<=tmp[1159]*kernel[0]+tmp[1160]*kernel[1]+tmp[1161]*kernel[2]+tmp[1259]*kernel[3]+tmp[1260]*kernel[4]+tmp[1261]*kernel[5]+tmp[1359]*kernel[6]+tmp[1360]*kernel[7]+tmp[1361]*kernel[8];
				ans[1261]<=tmp[1160]*kernel[0]+tmp[1161]*kernel[1]+tmp[1162]*kernel[2]+tmp[1260]*kernel[3]+tmp[1261]*kernel[4]+tmp[1262]*kernel[5]+tmp[1360]*kernel[6]+tmp[1361]*kernel[7]+tmp[1362]*kernel[8];
				ans[1262]<=tmp[1161]*kernel[0]+tmp[1162]*kernel[1]+tmp[1163]*kernel[2]+tmp[1261]*kernel[3]+tmp[1262]*kernel[4]+tmp[1263]*kernel[5]+tmp[1361]*kernel[6]+tmp[1362]*kernel[7]+tmp[1363]*kernel[8];
				ans[1263]<=tmp[1162]*kernel[0]+tmp[1163]*kernel[1]+tmp[1164]*kernel[2]+tmp[1262]*kernel[3]+tmp[1263]*kernel[4]+tmp[1264]*kernel[5]+tmp[1362]*kernel[6]+tmp[1363]*kernel[7]+tmp[1364]*kernel[8];
				ans[1264]<=tmp[1163]*kernel[0]+tmp[1164]*kernel[1]+tmp[1165]*kernel[2]+tmp[1263]*kernel[3]+tmp[1264]*kernel[4]+tmp[1265]*kernel[5]+tmp[1363]*kernel[6]+tmp[1364]*kernel[7]+tmp[1365]*kernel[8];
				ans[1265]<=tmp[1164]*kernel[0]+tmp[1165]*kernel[1]+tmp[1166]*kernel[2]+tmp[1264]*kernel[3]+tmp[1265]*kernel[4]+tmp[1266]*kernel[5]+tmp[1364]*kernel[6]+tmp[1365]*kernel[7]+tmp[1366]*kernel[8];
				ans[1266]<=tmp[1165]*kernel[0]+tmp[1166]*kernel[1]+tmp[1167]*kernel[2]+tmp[1265]*kernel[3]+tmp[1266]*kernel[4]+tmp[1267]*kernel[5]+tmp[1365]*kernel[6]+tmp[1366]*kernel[7]+tmp[1367]*kernel[8];
				ans[1267]<=tmp[1166]*kernel[0]+tmp[1167]*kernel[1]+tmp[1168]*kernel[2]+tmp[1266]*kernel[3]+tmp[1267]*kernel[4]+tmp[1268]*kernel[5]+tmp[1366]*kernel[6]+tmp[1367]*kernel[7]+tmp[1368]*kernel[8];
				ans[1268]<=tmp[1167]*kernel[0]+tmp[1168]*kernel[1]+tmp[1169]*kernel[2]+tmp[1267]*kernel[3]+tmp[1268]*kernel[4]+tmp[1269]*kernel[5]+tmp[1367]*kernel[6]+tmp[1368]*kernel[7]+tmp[1369]*kernel[8];
				ans[1269]<=tmp[1168]*kernel[0]+tmp[1169]*kernel[1]+tmp[1170]*kernel[2]+tmp[1268]*kernel[3]+tmp[1269]*kernel[4]+tmp[1270]*kernel[5]+tmp[1368]*kernel[6]+tmp[1369]*kernel[7]+tmp[1370]*kernel[8];
				ans[1270]<=tmp[1169]*kernel[0]+tmp[1170]*kernel[1]+tmp[1171]*kernel[2]+tmp[1269]*kernel[3]+tmp[1270]*kernel[4]+tmp[1271]*kernel[5]+tmp[1369]*kernel[6]+tmp[1370]*kernel[7]+tmp[1371]*kernel[8];
				ans[1271]<=tmp[1170]*kernel[0]+tmp[1171]*kernel[1]+tmp[1172]*kernel[2]+tmp[1270]*kernel[3]+tmp[1271]*kernel[4]+tmp[1272]*kernel[5]+tmp[1370]*kernel[6]+tmp[1371]*kernel[7]+tmp[1372]*kernel[8];
				ans[1272]<=tmp[1171]*kernel[0]+tmp[1172]*kernel[1]+tmp[1173]*kernel[2]+tmp[1271]*kernel[3]+tmp[1272]*kernel[4]+tmp[1273]*kernel[5]+tmp[1371]*kernel[6]+tmp[1372]*kernel[7]+tmp[1373]*kernel[8];
				ans[1273]<=tmp[1172]*kernel[0]+tmp[1173]*kernel[1]+tmp[1174]*kernel[2]+tmp[1272]*kernel[3]+tmp[1273]*kernel[4]+tmp[1274]*kernel[5]+tmp[1372]*kernel[6]+tmp[1373]*kernel[7]+tmp[1374]*kernel[8];
				ans[1274]<=tmp[1173]*kernel[0]+tmp[1174]*kernel[1]+tmp[1175]*kernel[2]+tmp[1273]*kernel[3]+tmp[1274]*kernel[4]+tmp[1275]*kernel[5]+tmp[1373]*kernel[6]+tmp[1374]*kernel[7]+tmp[1375]*kernel[8];
				ans[1275]<=tmp[1174]*kernel[0]+tmp[1175]*kernel[1]+tmp[1176]*kernel[2]+tmp[1274]*kernel[3]+tmp[1275]*kernel[4]+tmp[1276]*kernel[5]+tmp[1374]*kernel[6]+tmp[1375]*kernel[7]+tmp[1376]*kernel[8];
				ans[1276]<=tmp[1175]*kernel[0]+tmp[1176]*kernel[1]+tmp[1177]*kernel[2]+tmp[1275]*kernel[3]+tmp[1276]*kernel[4]+tmp[1277]*kernel[5]+tmp[1375]*kernel[6]+tmp[1376]*kernel[7]+tmp[1377]*kernel[8];
				ans[1277]<=tmp[1176]*kernel[0]+tmp[1177]*kernel[1]+tmp[1178]*kernel[2]+tmp[1276]*kernel[3]+tmp[1277]*kernel[4]+tmp[1278]*kernel[5]+tmp[1376]*kernel[6]+tmp[1377]*kernel[7]+tmp[1378]*kernel[8];
				ans[1278]<=tmp[1177]*kernel[0]+tmp[1178]*kernel[1]+tmp[1179]*kernel[2]+tmp[1277]*kernel[3]+tmp[1278]*kernel[4]+tmp[1279]*kernel[5]+tmp[1377]*kernel[6]+tmp[1378]*kernel[7]+tmp[1379]*kernel[8];
				ans[1279]<=tmp[1178]*kernel[0]+tmp[1179]*kernel[1]+tmp[1180]*kernel[2]+tmp[1278]*kernel[3]+tmp[1279]*kernel[4]+tmp[1280]*kernel[5]+tmp[1378]*kernel[6]+tmp[1379]*kernel[7]+tmp[1380]*kernel[8];
				ans[1280]<=tmp[1179]*kernel[0]+tmp[1180]*kernel[1]+tmp[1181]*kernel[2]+tmp[1279]*kernel[3]+tmp[1280]*kernel[4]+tmp[1281]*kernel[5]+tmp[1379]*kernel[6]+tmp[1380]*kernel[7]+tmp[1381]*kernel[8];
				ans[1281]<=tmp[1180]*kernel[0]+tmp[1181]*kernel[1]+tmp[1182]*kernel[2]+tmp[1280]*kernel[3]+tmp[1281]*kernel[4]+tmp[1282]*kernel[5]+tmp[1380]*kernel[6]+tmp[1381]*kernel[7]+tmp[1382]*kernel[8];
				ans[1282]<=tmp[1181]*kernel[0]+tmp[1182]*kernel[1]+tmp[1183]*kernel[2]+tmp[1281]*kernel[3]+tmp[1282]*kernel[4]+tmp[1283]*kernel[5]+tmp[1381]*kernel[6]+tmp[1382]*kernel[7]+tmp[1383]*kernel[8];
				ans[1283]<=tmp[1182]*kernel[0]+tmp[1183]*kernel[1]+tmp[1184]*kernel[2]+tmp[1282]*kernel[3]+tmp[1283]*kernel[4]+tmp[1284]*kernel[5]+tmp[1382]*kernel[6]+tmp[1383]*kernel[7]+tmp[1384]*kernel[8];
				ans[1284]<=tmp[1183]*kernel[0]+tmp[1184]*kernel[1]+tmp[1185]*kernel[2]+tmp[1283]*kernel[3]+tmp[1284]*kernel[4]+tmp[1285]*kernel[5]+tmp[1383]*kernel[6]+tmp[1384]*kernel[7]+tmp[1385]*kernel[8];
				ans[1285]<=tmp[1184]*kernel[0]+tmp[1185]*kernel[1]+tmp[1186]*kernel[2]+tmp[1284]*kernel[3]+tmp[1285]*kernel[4]+tmp[1286]*kernel[5]+tmp[1384]*kernel[6]+tmp[1385]*kernel[7]+tmp[1386]*kernel[8];
				ans[1286]<=tmp[1185]*kernel[0]+tmp[1186]*kernel[1]+tmp[1187]*kernel[2]+tmp[1285]*kernel[3]+tmp[1286]*kernel[4]+tmp[1287]*kernel[5]+tmp[1385]*kernel[6]+tmp[1386]*kernel[7]+tmp[1387]*kernel[8];
				ans[1287]<=tmp[1186]*kernel[0]+tmp[1187]*kernel[1]+tmp[1188]*kernel[2]+tmp[1286]*kernel[3]+tmp[1287]*kernel[4]+tmp[1288]*kernel[5]+tmp[1386]*kernel[6]+tmp[1387]*kernel[7]+tmp[1388]*kernel[8];
				ans[1288]<=tmp[1187]*kernel[0]+tmp[1188]*kernel[1]+tmp[1189]*kernel[2]+tmp[1287]*kernel[3]+tmp[1288]*kernel[4]+tmp[1289]*kernel[5]+tmp[1387]*kernel[6]+tmp[1388]*kernel[7]+tmp[1389]*kernel[8];
				ans[1289]<=tmp[1188]*kernel[0]+tmp[1189]*kernel[1]+tmp[1190]*kernel[2]+tmp[1288]*kernel[3]+tmp[1289]*kernel[4]+tmp[1290]*kernel[5]+tmp[1388]*kernel[6]+tmp[1389]*kernel[7]+tmp[1390]*kernel[8];
				ans[1290]<=tmp[1189]*kernel[0]+tmp[1190]*kernel[1]+tmp[1191]*kernel[2]+tmp[1289]*kernel[3]+tmp[1290]*kernel[4]+tmp[1291]*kernel[5]+tmp[1389]*kernel[6]+tmp[1390]*kernel[7]+tmp[1391]*kernel[8];
				ans[1291]<=tmp[1190]*kernel[0]+tmp[1191]*kernel[1]+tmp[1192]*kernel[2]+tmp[1290]*kernel[3]+tmp[1291]*kernel[4]+tmp[1292]*kernel[5]+tmp[1390]*kernel[6]+tmp[1391]*kernel[7]+tmp[1392]*kernel[8];
				ans[1292]<=tmp[1191]*kernel[0]+tmp[1192]*kernel[1]+tmp[1193]*kernel[2]+tmp[1291]*kernel[3]+tmp[1292]*kernel[4]+tmp[1293]*kernel[5]+tmp[1391]*kernel[6]+tmp[1392]*kernel[7]+tmp[1393]*kernel[8];
				ans[1293]<=tmp[1192]*kernel[0]+tmp[1193]*kernel[1]+tmp[1194]*kernel[2]+tmp[1292]*kernel[3]+tmp[1293]*kernel[4]+tmp[1294]*kernel[5]+tmp[1392]*kernel[6]+tmp[1393]*kernel[7]+tmp[1394]*kernel[8];
				ans[1294]<=tmp[1193]*kernel[0]+tmp[1194]*kernel[1]+tmp[1195]*kernel[2]+tmp[1293]*kernel[3]+tmp[1294]*kernel[4]+tmp[1295]*kernel[5]+tmp[1393]*kernel[6]+tmp[1394]*kernel[7]+tmp[1395]*kernel[8];
				ans[1295]<=tmp[1194]*kernel[0]+tmp[1195]*kernel[1]+tmp[1196]*kernel[2]+tmp[1294]*kernel[3]+tmp[1295]*kernel[4]+tmp[1296]*kernel[5]+tmp[1394]*kernel[6]+tmp[1395]*kernel[7]+tmp[1396]*kernel[8];
				ans[1296]<=tmp[1195]*kernel[0]+tmp[1196]*kernel[1]+tmp[1197]*kernel[2]+tmp[1295]*kernel[3]+tmp[1296]*kernel[4]+tmp[1297]*kernel[5]+tmp[1395]*kernel[6]+tmp[1396]*kernel[7]+tmp[1397]*kernel[8];
				ans[1297]<=tmp[1196]*kernel[0]+tmp[1197]*kernel[1]+tmp[1198]*kernel[2]+tmp[1296]*kernel[3]+tmp[1297]*kernel[4]+tmp[1298]*kernel[5]+tmp[1396]*kernel[6]+tmp[1397]*kernel[7]+tmp[1398]*kernel[8];
				ans[1298]<=tmp[1197]*kernel[0]+tmp[1198]*kernel[1]+tmp[1199]*kernel[2]+tmp[1297]*kernel[3]+tmp[1298]*kernel[4]+tmp[1299]*kernel[5]+tmp[1397]*kernel[6]+tmp[1398]*kernel[7]+tmp[1399]*kernel[8];
				ans[1299]<=tmp[1198]*kernel[0]+tmp[1199]*kernel[1]+tmp[1298]*kernel[3]+tmp[1299]*kernel[4]+tmp[1398]*kernel[6]+tmp[1399]*kernel[7];
				ans[1300]<=tmp[1200]*kernel[1]+tmp[1201]*kernel[2]+tmp[1300]*kernel[4]+tmp[1301]*kernel[5]+tmp[1400]*kernel[7]+tmp[1401]*kernel[8];
				ans[1301]<=tmp[1200]*kernel[0]+tmp[1201]*kernel[1]+tmp[1202]*kernel[2]+tmp[1300]*kernel[3]+tmp[1301]*kernel[4]+tmp[1302]*kernel[5]+tmp[1400]*kernel[6]+tmp[1401]*kernel[7]+tmp[1402]*kernel[8];
				ans[1302]<=tmp[1201]*kernel[0]+tmp[1202]*kernel[1]+tmp[1203]*kernel[2]+tmp[1301]*kernel[3]+tmp[1302]*kernel[4]+tmp[1303]*kernel[5]+tmp[1401]*kernel[6]+tmp[1402]*kernel[7]+tmp[1403]*kernel[8];
				ans[1303]<=tmp[1202]*kernel[0]+tmp[1203]*kernel[1]+tmp[1204]*kernel[2]+tmp[1302]*kernel[3]+tmp[1303]*kernel[4]+tmp[1304]*kernel[5]+tmp[1402]*kernel[6]+tmp[1403]*kernel[7]+tmp[1404]*kernel[8];
				ans[1304]<=tmp[1203]*kernel[0]+tmp[1204]*kernel[1]+tmp[1205]*kernel[2]+tmp[1303]*kernel[3]+tmp[1304]*kernel[4]+tmp[1305]*kernel[5]+tmp[1403]*kernel[6]+tmp[1404]*kernel[7]+tmp[1405]*kernel[8];
				ans[1305]<=tmp[1204]*kernel[0]+tmp[1205]*kernel[1]+tmp[1206]*kernel[2]+tmp[1304]*kernel[3]+tmp[1305]*kernel[4]+tmp[1306]*kernel[5]+tmp[1404]*kernel[6]+tmp[1405]*kernel[7]+tmp[1406]*kernel[8];
				ans[1306]<=tmp[1205]*kernel[0]+tmp[1206]*kernel[1]+tmp[1207]*kernel[2]+tmp[1305]*kernel[3]+tmp[1306]*kernel[4]+tmp[1307]*kernel[5]+tmp[1405]*kernel[6]+tmp[1406]*kernel[7]+tmp[1407]*kernel[8];
				ans[1307]<=tmp[1206]*kernel[0]+tmp[1207]*kernel[1]+tmp[1208]*kernel[2]+tmp[1306]*kernel[3]+tmp[1307]*kernel[4]+tmp[1308]*kernel[5]+tmp[1406]*kernel[6]+tmp[1407]*kernel[7]+tmp[1408]*kernel[8];
				ans[1308]<=tmp[1207]*kernel[0]+tmp[1208]*kernel[1]+tmp[1209]*kernel[2]+tmp[1307]*kernel[3]+tmp[1308]*kernel[4]+tmp[1309]*kernel[5]+tmp[1407]*kernel[6]+tmp[1408]*kernel[7]+tmp[1409]*kernel[8];
				ans[1309]<=tmp[1208]*kernel[0]+tmp[1209]*kernel[1]+tmp[1210]*kernel[2]+tmp[1308]*kernel[3]+tmp[1309]*kernel[4]+tmp[1310]*kernel[5]+tmp[1408]*kernel[6]+tmp[1409]*kernel[7]+tmp[1410]*kernel[8];
				ans[1310]<=tmp[1209]*kernel[0]+tmp[1210]*kernel[1]+tmp[1211]*kernel[2]+tmp[1309]*kernel[3]+tmp[1310]*kernel[4]+tmp[1311]*kernel[5]+tmp[1409]*kernel[6]+tmp[1410]*kernel[7]+tmp[1411]*kernel[8];
				ans[1311]<=tmp[1210]*kernel[0]+tmp[1211]*kernel[1]+tmp[1212]*kernel[2]+tmp[1310]*kernel[3]+tmp[1311]*kernel[4]+tmp[1312]*kernel[5]+tmp[1410]*kernel[6]+tmp[1411]*kernel[7]+tmp[1412]*kernel[8];
				ans[1312]<=tmp[1211]*kernel[0]+tmp[1212]*kernel[1]+tmp[1213]*kernel[2]+tmp[1311]*kernel[3]+tmp[1312]*kernel[4]+tmp[1313]*kernel[5]+tmp[1411]*kernel[6]+tmp[1412]*kernel[7]+tmp[1413]*kernel[8];
				ans[1313]<=tmp[1212]*kernel[0]+tmp[1213]*kernel[1]+tmp[1214]*kernel[2]+tmp[1312]*kernel[3]+tmp[1313]*kernel[4]+tmp[1314]*kernel[5]+tmp[1412]*kernel[6]+tmp[1413]*kernel[7]+tmp[1414]*kernel[8];
				ans[1314]<=tmp[1213]*kernel[0]+tmp[1214]*kernel[1]+tmp[1215]*kernel[2]+tmp[1313]*kernel[3]+tmp[1314]*kernel[4]+tmp[1315]*kernel[5]+tmp[1413]*kernel[6]+tmp[1414]*kernel[7]+tmp[1415]*kernel[8];
				ans[1315]<=tmp[1214]*kernel[0]+tmp[1215]*kernel[1]+tmp[1216]*kernel[2]+tmp[1314]*kernel[3]+tmp[1315]*kernel[4]+tmp[1316]*kernel[5]+tmp[1414]*kernel[6]+tmp[1415]*kernel[7]+tmp[1416]*kernel[8];
				ans[1316]<=tmp[1215]*kernel[0]+tmp[1216]*kernel[1]+tmp[1217]*kernel[2]+tmp[1315]*kernel[3]+tmp[1316]*kernel[4]+tmp[1317]*kernel[5]+tmp[1415]*kernel[6]+tmp[1416]*kernel[7]+tmp[1417]*kernel[8];
				ans[1317]<=tmp[1216]*kernel[0]+tmp[1217]*kernel[1]+tmp[1218]*kernel[2]+tmp[1316]*kernel[3]+tmp[1317]*kernel[4]+tmp[1318]*kernel[5]+tmp[1416]*kernel[6]+tmp[1417]*kernel[7]+tmp[1418]*kernel[8];
				ans[1318]<=tmp[1217]*kernel[0]+tmp[1218]*kernel[1]+tmp[1219]*kernel[2]+tmp[1317]*kernel[3]+tmp[1318]*kernel[4]+tmp[1319]*kernel[5]+tmp[1417]*kernel[6]+tmp[1418]*kernel[7]+tmp[1419]*kernel[8];
				ans[1319]<=tmp[1218]*kernel[0]+tmp[1219]*kernel[1]+tmp[1220]*kernel[2]+tmp[1318]*kernel[3]+tmp[1319]*kernel[4]+tmp[1320]*kernel[5]+tmp[1418]*kernel[6]+tmp[1419]*kernel[7]+tmp[1420]*kernel[8];
				ans[1320]<=tmp[1219]*kernel[0]+tmp[1220]*kernel[1]+tmp[1221]*kernel[2]+tmp[1319]*kernel[3]+tmp[1320]*kernel[4]+tmp[1321]*kernel[5]+tmp[1419]*kernel[6]+tmp[1420]*kernel[7]+tmp[1421]*kernel[8];
				ans[1321]<=tmp[1220]*kernel[0]+tmp[1221]*kernel[1]+tmp[1222]*kernel[2]+tmp[1320]*kernel[3]+tmp[1321]*kernel[4]+tmp[1322]*kernel[5]+tmp[1420]*kernel[6]+tmp[1421]*kernel[7]+tmp[1422]*kernel[8];
				ans[1322]<=tmp[1221]*kernel[0]+tmp[1222]*kernel[1]+tmp[1223]*kernel[2]+tmp[1321]*kernel[3]+tmp[1322]*kernel[4]+tmp[1323]*kernel[5]+tmp[1421]*kernel[6]+tmp[1422]*kernel[7]+tmp[1423]*kernel[8];
				ans[1323]<=tmp[1222]*kernel[0]+tmp[1223]*kernel[1]+tmp[1224]*kernel[2]+tmp[1322]*kernel[3]+tmp[1323]*kernel[4]+tmp[1324]*kernel[5]+tmp[1422]*kernel[6]+tmp[1423]*kernel[7]+tmp[1424]*kernel[8];
				ans[1324]<=tmp[1223]*kernel[0]+tmp[1224]*kernel[1]+tmp[1225]*kernel[2]+tmp[1323]*kernel[3]+tmp[1324]*kernel[4]+tmp[1325]*kernel[5]+tmp[1423]*kernel[6]+tmp[1424]*kernel[7]+tmp[1425]*kernel[8];
				ans[1325]<=tmp[1224]*kernel[0]+tmp[1225]*kernel[1]+tmp[1226]*kernel[2]+tmp[1324]*kernel[3]+tmp[1325]*kernel[4]+tmp[1326]*kernel[5]+tmp[1424]*kernel[6]+tmp[1425]*kernel[7]+tmp[1426]*kernel[8];
				ans[1326]<=tmp[1225]*kernel[0]+tmp[1226]*kernel[1]+tmp[1227]*kernel[2]+tmp[1325]*kernel[3]+tmp[1326]*kernel[4]+tmp[1327]*kernel[5]+tmp[1425]*kernel[6]+tmp[1426]*kernel[7]+tmp[1427]*kernel[8];
				ans[1327]<=tmp[1226]*kernel[0]+tmp[1227]*kernel[1]+tmp[1228]*kernel[2]+tmp[1326]*kernel[3]+tmp[1327]*kernel[4]+tmp[1328]*kernel[5]+tmp[1426]*kernel[6]+tmp[1427]*kernel[7]+tmp[1428]*kernel[8];
				ans[1328]<=tmp[1227]*kernel[0]+tmp[1228]*kernel[1]+tmp[1229]*kernel[2]+tmp[1327]*kernel[3]+tmp[1328]*kernel[4]+tmp[1329]*kernel[5]+tmp[1427]*kernel[6]+tmp[1428]*kernel[7]+tmp[1429]*kernel[8];
				ans[1329]<=tmp[1228]*kernel[0]+tmp[1229]*kernel[1]+tmp[1230]*kernel[2]+tmp[1328]*kernel[3]+tmp[1329]*kernel[4]+tmp[1330]*kernel[5]+tmp[1428]*kernel[6]+tmp[1429]*kernel[7]+tmp[1430]*kernel[8];
				ans[1330]<=tmp[1229]*kernel[0]+tmp[1230]*kernel[1]+tmp[1231]*kernel[2]+tmp[1329]*kernel[3]+tmp[1330]*kernel[4]+tmp[1331]*kernel[5]+tmp[1429]*kernel[6]+tmp[1430]*kernel[7]+tmp[1431]*kernel[8];
				ans[1331]<=tmp[1230]*kernel[0]+tmp[1231]*kernel[1]+tmp[1232]*kernel[2]+tmp[1330]*kernel[3]+tmp[1331]*kernel[4]+tmp[1332]*kernel[5]+tmp[1430]*kernel[6]+tmp[1431]*kernel[7]+tmp[1432]*kernel[8];
				ans[1332]<=tmp[1231]*kernel[0]+tmp[1232]*kernel[1]+tmp[1233]*kernel[2]+tmp[1331]*kernel[3]+tmp[1332]*kernel[4]+tmp[1333]*kernel[5]+tmp[1431]*kernel[6]+tmp[1432]*kernel[7]+tmp[1433]*kernel[8];
				ans[1333]<=tmp[1232]*kernel[0]+tmp[1233]*kernel[1]+tmp[1234]*kernel[2]+tmp[1332]*kernel[3]+tmp[1333]*kernel[4]+tmp[1334]*kernel[5]+tmp[1432]*kernel[6]+tmp[1433]*kernel[7]+tmp[1434]*kernel[8];
				ans[1334]<=tmp[1233]*kernel[0]+tmp[1234]*kernel[1]+tmp[1235]*kernel[2]+tmp[1333]*kernel[3]+tmp[1334]*kernel[4]+tmp[1335]*kernel[5]+tmp[1433]*kernel[6]+tmp[1434]*kernel[7]+tmp[1435]*kernel[8];
				ans[1335]<=tmp[1234]*kernel[0]+tmp[1235]*kernel[1]+tmp[1236]*kernel[2]+tmp[1334]*kernel[3]+tmp[1335]*kernel[4]+tmp[1336]*kernel[5]+tmp[1434]*kernel[6]+tmp[1435]*kernel[7]+tmp[1436]*kernel[8];
				ans[1336]<=tmp[1235]*kernel[0]+tmp[1236]*kernel[1]+tmp[1237]*kernel[2]+tmp[1335]*kernel[3]+tmp[1336]*kernel[4]+tmp[1337]*kernel[5]+tmp[1435]*kernel[6]+tmp[1436]*kernel[7]+tmp[1437]*kernel[8];
				ans[1337]<=tmp[1236]*kernel[0]+tmp[1237]*kernel[1]+tmp[1238]*kernel[2]+tmp[1336]*kernel[3]+tmp[1337]*kernel[4]+tmp[1338]*kernel[5]+tmp[1436]*kernel[6]+tmp[1437]*kernel[7]+tmp[1438]*kernel[8];
				ans[1338]<=tmp[1237]*kernel[0]+tmp[1238]*kernel[1]+tmp[1239]*kernel[2]+tmp[1337]*kernel[3]+tmp[1338]*kernel[4]+tmp[1339]*kernel[5]+tmp[1437]*kernel[6]+tmp[1438]*kernel[7]+tmp[1439]*kernel[8];
				ans[1339]<=tmp[1238]*kernel[0]+tmp[1239]*kernel[1]+tmp[1240]*kernel[2]+tmp[1338]*kernel[3]+tmp[1339]*kernel[4]+tmp[1340]*kernel[5]+tmp[1438]*kernel[6]+tmp[1439]*kernel[7]+tmp[1440]*kernel[8];
				ans[1340]<=tmp[1239]*kernel[0]+tmp[1240]*kernel[1]+tmp[1241]*kernel[2]+tmp[1339]*kernel[3]+tmp[1340]*kernel[4]+tmp[1341]*kernel[5]+tmp[1439]*kernel[6]+tmp[1440]*kernel[7]+tmp[1441]*kernel[8];
				ans[1341]<=tmp[1240]*kernel[0]+tmp[1241]*kernel[1]+tmp[1242]*kernel[2]+tmp[1340]*kernel[3]+tmp[1341]*kernel[4]+tmp[1342]*kernel[5]+tmp[1440]*kernel[6]+tmp[1441]*kernel[7]+tmp[1442]*kernel[8];
				ans[1342]<=tmp[1241]*kernel[0]+tmp[1242]*kernel[1]+tmp[1243]*kernel[2]+tmp[1341]*kernel[3]+tmp[1342]*kernel[4]+tmp[1343]*kernel[5]+tmp[1441]*kernel[6]+tmp[1442]*kernel[7]+tmp[1443]*kernel[8];
				ans[1343]<=tmp[1242]*kernel[0]+tmp[1243]*kernel[1]+tmp[1244]*kernel[2]+tmp[1342]*kernel[3]+tmp[1343]*kernel[4]+tmp[1344]*kernel[5]+tmp[1442]*kernel[6]+tmp[1443]*kernel[7]+tmp[1444]*kernel[8];
				ans[1344]<=tmp[1243]*kernel[0]+tmp[1244]*kernel[1]+tmp[1245]*kernel[2]+tmp[1343]*kernel[3]+tmp[1344]*kernel[4]+tmp[1345]*kernel[5]+tmp[1443]*kernel[6]+tmp[1444]*kernel[7]+tmp[1445]*kernel[8];
				ans[1345]<=tmp[1244]*kernel[0]+tmp[1245]*kernel[1]+tmp[1246]*kernel[2]+tmp[1344]*kernel[3]+tmp[1345]*kernel[4]+tmp[1346]*kernel[5]+tmp[1444]*kernel[6]+tmp[1445]*kernel[7]+tmp[1446]*kernel[8];
				ans[1346]<=tmp[1245]*kernel[0]+tmp[1246]*kernel[1]+tmp[1247]*kernel[2]+tmp[1345]*kernel[3]+tmp[1346]*kernel[4]+tmp[1347]*kernel[5]+tmp[1445]*kernel[6]+tmp[1446]*kernel[7]+tmp[1447]*kernel[8];
				ans[1347]<=tmp[1246]*kernel[0]+tmp[1247]*kernel[1]+tmp[1248]*kernel[2]+tmp[1346]*kernel[3]+tmp[1347]*kernel[4]+tmp[1348]*kernel[5]+tmp[1446]*kernel[6]+tmp[1447]*kernel[7]+tmp[1448]*kernel[8];
				ans[1348]<=tmp[1247]*kernel[0]+tmp[1248]*kernel[1]+tmp[1249]*kernel[2]+tmp[1347]*kernel[3]+tmp[1348]*kernel[4]+tmp[1349]*kernel[5]+tmp[1447]*kernel[6]+tmp[1448]*kernel[7]+tmp[1449]*kernel[8];
				ans[1349]<=tmp[1248]*kernel[0]+tmp[1249]*kernel[1]+tmp[1250]*kernel[2]+tmp[1348]*kernel[3]+tmp[1349]*kernel[4]+tmp[1350]*kernel[5]+tmp[1448]*kernel[6]+tmp[1449]*kernel[7]+tmp[1450]*kernel[8];
				ans[1350]<=tmp[1249]*kernel[0]+tmp[1250]*kernel[1]+tmp[1251]*kernel[2]+tmp[1349]*kernel[3]+tmp[1350]*kernel[4]+tmp[1351]*kernel[5]+tmp[1449]*kernel[6]+tmp[1450]*kernel[7]+tmp[1451]*kernel[8];
				ans[1351]<=tmp[1250]*kernel[0]+tmp[1251]*kernel[1]+tmp[1252]*kernel[2]+tmp[1350]*kernel[3]+tmp[1351]*kernel[4]+tmp[1352]*kernel[5]+tmp[1450]*kernel[6]+tmp[1451]*kernel[7]+tmp[1452]*kernel[8];
				ans[1352]<=tmp[1251]*kernel[0]+tmp[1252]*kernel[1]+tmp[1253]*kernel[2]+tmp[1351]*kernel[3]+tmp[1352]*kernel[4]+tmp[1353]*kernel[5]+tmp[1451]*kernel[6]+tmp[1452]*kernel[7]+tmp[1453]*kernel[8];
				ans[1353]<=tmp[1252]*kernel[0]+tmp[1253]*kernel[1]+tmp[1254]*kernel[2]+tmp[1352]*kernel[3]+tmp[1353]*kernel[4]+tmp[1354]*kernel[5]+tmp[1452]*kernel[6]+tmp[1453]*kernel[7]+tmp[1454]*kernel[8];
				ans[1354]<=tmp[1253]*kernel[0]+tmp[1254]*kernel[1]+tmp[1255]*kernel[2]+tmp[1353]*kernel[3]+tmp[1354]*kernel[4]+tmp[1355]*kernel[5]+tmp[1453]*kernel[6]+tmp[1454]*kernel[7]+tmp[1455]*kernel[8];
				ans[1355]<=tmp[1254]*kernel[0]+tmp[1255]*kernel[1]+tmp[1256]*kernel[2]+tmp[1354]*kernel[3]+tmp[1355]*kernel[4]+tmp[1356]*kernel[5]+tmp[1454]*kernel[6]+tmp[1455]*kernel[7]+tmp[1456]*kernel[8];
				ans[1356]<=tmp[1255]*kernel[0]+tmp[1256]*kernel[1]+tmp[1257]*kernel[2]+tmp[1355]*kernel[3]+tmp[1356]*kernel[4]+tmp[1357]*kernel[5]+tmp[1455]*kernel[6]+tmp[1456]*kernel[7]+tmp[1457]*kernel[8];
				ans[1357]<=tmp[1256]*kernel[0]+tmp[1257]*kernel[1]+tmp[1258]*kernel[2]+tmp[1356]*kernel[3]+tmp[1357]*kernel[4]+tmp[1358]*kernel[5]+tmp[1456]*kernel[6]+tmp[1457]*kernel[7]+tmp[1458]*kernel[8];
				ans[1358]<=tmp[1257]*kernel[0]+tmp[1258]*kernel[1]+tmp[1259]*kernel[2]+tmp[1357]*kernel[3]+tmp[1358]*kernel[4]+tmp[1359]*kernel[5]+tmp[1457]*kernel[6]+tmp[1458]*kernel[7]+tmp[1459]*kernel[8];
				ans[1359]<=tmp[1258]*kernel[0]+tmp[1259]*kernel[1]+tmp[1260]*kernel[2]+tmp[1358]*kernel[3]+tmp[1359]*kernel[4]+tmp[1360]*kernel[5]+tmp[1458]*kernel[6]+tmp[1459]*kernel[7]+tmp[1460]*kernel[8];
				ans[1360]<=tmp[1259]*kernel[0]+tmp[1260]*kernel[1]+tmp[1261]*kernel[2]+tmp[1359]*kernel[3]+tmp[1360]*kernel[4]+tmp[1361]*kernel[5]+tmp[1459]*kernel[6]+tmp[1460]*kernel[7]+tmp[1461]*kernel[8];
				ans[1361]<=tmp[1260]*kernel[0]+tmp[1261]*kernel[1]+tmp[1262]*kernel[2]+tmp[1360]*kernel[3]+tmp[1361]*kernel[4]+tmp[1362]*kernel[5]+tmp[1460]*kernel[6]+tmp[1461]*kernel[7]+tmp[1462]*kernel[8];
				ans[1362]<=tmp[1261]*kernel[0]+tmp[1262]*kernel[1]+tmp[1263]*kernel[2]+tmp[1361]*kernel[3]+tmp[1362]*kernel[4]+tmp[1363]*kernel[5]+tmp[1461]*kernel[6]+tmp[1462]*kernel[7]+tmp[1463]*kernel[8];
				ans[1363]<=tmp[1262]*kernel[0]+tmp[1263]*kernel[1]+tmp[1264]*kernel[2]+tmp[1362]*kernel[3]+tmp[1363]*kernel[4]+tmp[1364]*kernel[5]+tmp[1462]*kernel[6]+tmp[1463]*kernel[7]+tmp[1464]*kernel[8];
				ans[1364]<=tmp[1263]*kernel[0]+tmp[1264]*kernel[1]+tmp[1265]*kernel[2]+tmp[1363]*kernel[3]+tmp[1364]*kernel[4]+tmp[1365]*kernel[5]+tmp[1463]*kernel[6]+tmp[1464]*kernel[7]+tmp[1465]*kernel[8];
				ans[1365]<=tmp[1264]*kernel[0]+tmp[1265]*kernel[1]+tmp[1266]*kernel[2]+tmp[1364]*kernel[3]+tmp[1365]*kernel[4]+tmp[1366]*kernel[5]+tmp[1464]*kernel[6]+tmp[1465]*kernel[7]+tmp[1466]*kernel[8];
				ans[1366]<=tmp[1265]*kernel[0]+tmp[1266]*kernel[1]+tmp[1267]*kernel[2]+tmp[1365]*kernel[3]+tmp[1366]*kernel[4]+tmp[1367]*kernel[5]+tmp[1465]*kernel[6]+tmp[1466]*kernel[7]+tmp[1467]*kernel[8];
				ans[1367]<=tmp[1266]*kernel[0]+tmp[1267]*kernel[1]+tmp[1268]*kernel[2]+tmp[1366]*kernel[3]+tmp[1367]*kernel[4]+tmp[1368]*kernel[5]+tmp[1466]*kernel[6]+tmp[1467]*kernel[7]+tmp[1468]*kernel[8];
				ans[1368]<=tmp[1267]*kernel[0]+tmp[1268]*kernel[1]+tmp[1269]*kernel[2]+tmp[1367]*kernel[3]+tmp[1368]*kernel[4]+tmp[1369]*kernel[5]+tmp[1467]*kernel[6]+tmp[1468]*kernel[7]+tmp[1469]*kernel[8];
				ans[1369]<=tmp[1268]*kernel[0]+tmp[1269]*kernel[1]+tmp[1270]*kernel[2]+tmp[1368]*kernel[3]+tmp[1369]*kernel[4]+tmp[1370]*kernel[5]+tmp[1468]*kernel[6]+tmp[1469]*kernel[7]+tmp[1470]*kernel[8];
				ans[1370]<=tmp[1269]*kernel[0]+tmp[1270]*kernel[1]+tmp[1271]*kernel[2]+tmp[1369]*kernel[3]+tmp[1370]*kernel[4]+tmp[1371]*kernel[5]+tmp[1469]*kernel[6]+tmp[1470]*kernel[7]+tmp[1471]*kernel[8];
				ans[1371]<=tmp[1270]*kernel[0]+tmp[1271]*kernel[1]+tmp[1272]*kernel[2]+tmp[1370]*kernel[3]+tmp[1371]*kernel[4]+tmp[1372]*kernel[5]+tmp[1470]*kernel[6]+tmp[1471]*kernel[7]+tmp[1472]*kernel[8];
				ans[1372]<=tmp[1271]*kernel[0]+tmp[1272]*kernel[1]+tmp[1273]*kernel[2]+tmp[1371]*kernel[3]+tmp[1372]*kernel[4]+tmp[1373]*kernel[5]+tmp[1471]*kernel[6]+tmp[1472]*kernel[7]+tmp[1473]*kernel[8];
				ans[1373]<=tmp[1272]*kernel[0]+tmp[1273]*kernel[1]+tmp[1274]*kernel[2]+tmp[1372]*kernel[3]+tmp[1373]*kernel[4]+tmp[1374]*kernel[5]+tmp[1472]*kernel[6]+tmp[1473]*kernel[7]+tmp[1474]*kernel[8];
				ans[1374]<=tmp[1273]*kernel[0]+tmp[1274]*kernel[1]+tmp[1275]*kernel[2]+tmp[1373]*kernel[3]+tmp[1374]*kernel[4]+tmp[1375]*kernel[5]+tmp[1473]*kernel[6]+tmp[1474]*kernel[7]+tmp[1475]*kernel[8];
				ans[1375]<=tmp[1274]*kernel[0]+tmp[1275]*kernel[1]+tmp[1276]*kernel[2]+tmp[1374]*kernel[3]+tmp[1375]*kernel[4]+tmp[1376]*kernel[5]+tmp[1474]*kernel[6]+tmp[1475]*kernel[7]+tmp[1476]*kernel[8];
				ans[1376]<=tmp[1275]*kernel[0]+tmp[1276]*kernel[1]+tmp[1277]*kernel[2]+tmp[1375]*kernel[3]+tmp[1376]*kernel[4]+tmp[1377]*kernel[5]+tmp[1475]*kernel[6]+tmp[1476]*kernel[7]+tmp[1477]*kernel[8];
				ans[1377]<=tmp[1276]*kernel[0]+tmp[1277]*kernel[1]+tmp[1278]*kernel[2]+tmp[1376]*kernel[3]+tmp[1377]*kernel[4]+tmp[1378]*kernel[5]+tmp[1476]*kernel[6]+tmp[1477]*kernel[7]+tmp[1478]*kernel[8];
				ans[1378]<=tmp[1277]*kernel[0]+tmp[1278]*kernel[1]+tmp[1279]*kernel[2]+tmp[1377]*kernel[3]+tmp[1378]*kernel[4]+tmp[1379]*kernel[5]+tmp[1477]*kernel[6]+tmp[1478]*kernel[7]+tmp[1479]*kernel[8];
				ans[1379]<=tmp[1278]*kernel[0]+tmp[1279]*kernel[1]+tmp[1280]*kernel[2]+tmp[1378]*kernel[3]+tmp[1379]*kernel[4]+tmp[1380]*kernel[5]+tmp[1478]*kernel[6]+tmp[1479]*kernel[7]+tmp[1480]*kernel[8];
				ans[1380]<=tmp[1279]*kernel[0]+tmp[1280]*kernel[1]+tmp[1281]*kernel[2]+tmp[1379]*kernel[3]+tmp[1380]*kernel[4]+tmp[1381]*kernel[5]+tmp[1479]*kernel[6]+tmp[1480]*kernel[7]+tmp[1481]*kernel[8];
				ans[1381]<=tmp[1280]*kernel[0]+tmp[1281]*kernel[1]+tmp[1282]*kernel[2]+tmp[1380]*kernel[3]+tmp[1381]*kernel[4]+tmp[1382]*kernel[5]+tmp[1480]*kernel[6]+tmp[1481]*kernel[7]+tmp[1482]*kernel[8];
				ans[1382]<=tmp[1281]*kernel[0]+tmp[1282]*kernel[1]+tmp[1283]*kernel[2]+tmp[1381]*kernel[3]+tmp[1382]*kernel[4]+tmp[1383]*kernel[5]+tmp[1481]*kernel[6]+tmp[1482]*kernel[7]+tmp[1483]*kernel[8];
				ans[1383]<=tmp[1282]*kernel[0]+tmp[1283]*kernel[1]+tmp[1284]*kernel[2]+tmp[1382]*kernel[3]+tmp[1383]*kernel[4]+tmp[1384]*kernel[5]+tmp[1482]*kernel[6]+tmp[1483]*kernel[7]+tmp[1484]*kernel[8];
				ans[1384]<=tmp[1283]*kernel[0]+tmp[1284]*kernel[1]+tmp[1285]*kernel[2]+tmp[1383]*kernel[3]+tmp[1384]*kernel[4]+tmp[1385]*kernel[5]+tmp[1483]*kernel[6]+tmp[1484]*kernel[7]+tmp[1485]*kernel[8];
				ans[1385]<=tmp[1284]*kernel[0]+tmp[1285]*kernel[1]+tmp[1286]*kernel[2]+tmp[1384]*kernel[3]+tmp[1385]*kernel[4]+tmp[1386]*kernel[5]+tmp[1484]*kernel[6]+tmp[1485]*kernel[7]+tmp[1486]*kernel[8];
				ans[1386]<=tmp[1285]*kernel[0]+tmp[1286]*kernel[1]+tmp[1287]*kernel[2]+tmp[1385]*kernel[3]+tmp[1386]*kernel[4]+tmp[1387]*kernel[5]+tmp[1485]*kernel[6]+tmp[1486]*kernel[7]+tmp[1487]*kernel[8];
				ans[1387]<=tmp[1286]*kernel[0]+tmp[1287]*kernel[1]+tmp[1288]*kernel[2]+tmp[1386]*kernel[3]+tmp[1387]*kernel[4]+tmp[1388]*kernel[5]+tmp[1486]*kernel[6]+tmp[1487]*kernel[7]+tmp[1488]*kernel[8];
				ans[1388]<=tmp[1287]*kernel[0]+tmp[1288]*kernel[1]+tmp[1289]*kernel[2]+tmp[1387]*kernel[3]+tmp[1388]*kernel[4]+tmp[1389]*kernel[5]+tmp[1487]*kernel[6]+tmp[1488]*kernel[7]+tmp[1489]*kernel[8];
				ans[1389]<=tmp[1288]*kernel[0]+tmp[1289]*kernel[1]+tmp[1290]*kernel[2]+tmp[1388]*kernel[3]+tmp[1389]*kernel[4]+tmp[1390]*kernel[5]+tmp[1488]*kernel[6]+tmp[1489]*kernel[7]+tmp[1490]*kernel[8];
				ans[1390]<=tmp[1289]*kernel[0]+tmp[1290]*kernel[1]+tmp[1291]*kernel[2]+tmp[1389]*kernel[3]+tmp[1390]*kernel[4]+tmp[1391]*kernel[5]+tmp[1489]*kernel[6]+tmp[1490]*kernel[7]+tmp[1491]*kernel[8];
				ans[1391]<=tmp[1290]*kernel[0]+tmp[1291]*kernel[1]+tmp[1292]*kernel[2]+tmp[1390]*kernel[3]+tmp[1391]*kernel[4]+tmp[1392]*kernel[5]+tmp[1490]*kernel[6]+tmp[1491]*kernel[7]+tmp[1492]*kernel[8];
				ans[1392]<=tmp[1291]*kernel[0]+tmp[1292]*kernel[1]+tmp[1293]*kernel[2]+tmp[1391]*kernel[3]+tmp[1392]*kernel[4]+tmp[1393]*kernel[5]+tmp[1491]*kernel[6]+tmp[1492]*kernel[7]+tmp[1493]*kernel[8];
				ans[1393]<=tmp[1292]*kernel[0]+tmp[1293]*kernel[1]+tmp[1294]*kernel[2]+tmp[1392]*kernel[3]+tmp[1393]*kernel[4]+tmp[1394]*kernel[5]+tmp[1492]*kernel[6]+tmp[1493]*kernel[7]+tmp[1494]*kernel[8];
				ans[1394]<=tmp[1293]*kernel[0]+tmp[1294]*kernel[1]+tmp[1295]*kernel[2]+tmp[1393]*kernel[3]+tmp[1394]*kernel[4]+tmp[1395]*kernel[5]+tmp[1493]*kernel[6]+tmp[1494]*kernel[7]+tmp[1495]*kernel[8];
				ans[1395]<=tmp[1294]*kernel[0]+tmp[1295]*kernel[1]+tmp[1296]*kernel[2]+tmp[1394]*kernel[3]+tmp[1395]*kernel[4]+tmp[1396]*kernel[5]+tmp[1494]*kernel[6]+tmp[1495]*kernel[7]+tmp[1496]*kernel[8];
				ans[1396]<=tmp[1295]*kernel[0]+tmp[1296]*kernel[1]+tmp[1297]*kernel[2]+tmp[1395]*kernel[3]+tmp[1396]*kernel[4]+tmp[1397]*kernel[5]+tmp[1495]*kernel[6]+tmp[1496]*kernel[7]+tmp[1497]*kernel[8];
				ans[1397]<=tmp[1296]*kernel[0]+tmp[1297]*kernel[1]+tmp[1298]*kernel[2]+tmp[1396]*kernel[3]+tmp[1397]*kernel[4]+tmp[1398]*kernel[5]+tmp[1496]*kernel[6]+tmp[1497]*kernel[7]+tmp[1498]*kernel[8];
				ans[1398]<=tmp[1297]*kernel[0]+tmp[1298]*kernel[1]+tmp[1299]*kernel[2]+tmp[1397]*kernel[3]+tmp[1398]*kernel[4]+tmp[1399]*kernel[5]+tmp[1497]*kernel[6]+tmp[1498]*kernel[7]+tmp[1499]*kernel[8];
				ans[1399]<=tmp[1298]*kernel[0]+tmp[1299]*kernel[1]+tmp[1398]*kernel[3]+tmp[1399]*kernel[4]+tmp[1498]*kernel[6]+tmp[1499]*kernel[7];
				ans[1400]<=tmp[1300]*kernel[1]+tmp[1301]*kernel[2]+tmp[1400]*kernel[4]+tmp[1401]*kernel[5]+tmp[1500]*kernel[7]+tmp[1501]*kernel[8];
				ans[1401]<=tmp[1300]*kernel[0]+tmp[1301]*kernel[1]+tmp[1302]*kernel[2]+tmp[1400]*kernel[3]+tmp[1401]*kernel[4]+tmp[1402]*kernel[5]+tmp[1500]*kernel[6]+tmp[1501]*kernel[7]+tmp[1502]*kernel[8];
				ans[1402]<=tmp[1301]*kernel[0]+tmp[1302]*kernel[1]+tmp[1303]*kernel[2]+tmp[1401]*kernel[3]+tmp[1402]*kernel[4]+tmp[1403]*kernel[5]+tmp[1501]*kernel[6]+tmp[1502]*kernel[7]+tmp[1503]*kernel[8];
				ans[1403]<=tmp[1302]*kernel[0]+tmp[1303]*kernel[1]+tmp[1304]*kernel[2]+tmp[1402]*kernel[3]+tmp[1403]*kernel[4]+tmp[1404]*kernel[5]+tmp[1502]*kernel[6]+tmp[1503]*kernel[7]+tmp[1504]*kernel[8];
				ans[1404]<=tmp[1303]*kernel[0]+tmp[1304]*kernel[1]+tmp[1305]*kernel[2]+tmp[1403]*kernel[3]+tmp[1404]*kernel[4]+tmp[1405]*kernel[5]+tmp[1503]*kernel[6]+tmp[1504]*kernel[7]+tmp[1505]*kernel[8];
				ans[1405]<=tmp[1304]*kernel[0]+tmp[1305]*kernel[1]+tmp[1306]*kernel[2]+tmp[1404]*kernel[3]+tmp[1405]*kernel[4]+tmp[1406]*kernel[5]+tmp[1504]*kernel[6]+tmp[1505]*kernel[7]+tmp[1506]*kernel[8];
				ans[1406]<=tmp[1305]*kernel[0]+tmp[1306]*kernel[1]+tmp[1307]*kernel[2]+tmp[1405]*kernel[3]+tmp[1406]*kernel[4]+tmp[1407]*kernel[5]+tmp[1505]*kernel[6]+tmp[1506]*kernel[7]+tmp[1507]*kernel[8];
				ans[1407]<=tmp[1306]*kernel[0]+tmp[1307]*kernel[1]+tmp[1308]*kernel[2]+tmp[1406]*kernel[3]+tmp[1407]*kernel[4]+tmp[1408]*kernel[5]+tmp[1506]*kernel[6]+tmp[1507]*kernel[7]+tmp[1508]*kernel[8];
				ans[1408]<=tmp[1307]*kernel[0]+tmp[1308]*kernel[1]+tmp[1309]*kernel[2]+tmp[1407]*kernel[3]+tmp[1408]*kernel[4]+tmp[1409]*kernel[5]+tmp[1507]*kernel[6]+tmp[1508]*kernel[7]+tmp[1509]*kernel[8];
				ans[1409]<=tmp[1308]*kernel[0]+tmp[1309]*kernel[1]+tmp[1310]*kernel[2]+tmp[1408]*kernel[3]+tmp[1409]*kernel[4]+tmp[1410]*kernel[5]+tmp[1508]*kernel[6]+tmp[1509]*kernel[7]+tmp[1510]*kernel[8];
				ans[1410]<=tmp[1309]*kernel[0]+tmp[1310]*kernel[1]+tmp[1311]*kernel[2]+tmp[1409]*kernel[3]+tmp[1410]*kernel[4]+tmp[1411]*kernel[5]+tmp[1509]*kernel[6]+tmp[1510]*kernel[7]+tmp[1511]*kernel[8];
				ans[1411]<=tmp[1310]*kernel[0]+tmp[1311]*kernel[1]+tmp[1312]*kernel[2]+tmp[1410]*kernel[3]+tmp[1411]*kernel[4]+tmp[1412]*kernel[5]+tmp[1510]*kernel[6]+tmp[1511]*kernel[7]+tmp[1512]*kernel[8];
				ans[1412]<=tmp[1311]*kernel[0]+tmp[1312]*kernel[1]+tmp[1313]*kernel[2]+tmp[1411]*kernel[3]+tmp[1412]*kernel[4]+tmp[1413]*kernel[5]+tmp[1511]*kernel[6]+tmp[1512]*kernel[7]+tmp[1513]*kernel[8];
				ans[1413]<=tmp[1312]*kernel[0]+tmp[1313]*kernel[1]+tmp[1314]*kernel[2]+tmp[1412]*kernel[3]+tmp[1413]*kernel[4]+tmp[1414]*kernel[5]+tmp[1512]*kernel[6]+tmp[1513]*kernel[7]+tmp[1514]*kernel[8];
				ans[1414]<=tmp[1313]*kernel[0]+tmp[1314]*kernel[1]+tmp[1315]*kernel[2]+tmp[1413]*kernel[3]+tmp[1414]*kernel[4]+tmp[1415]*kernel[5]+tmp[1513]*kernel[6]+tmp[1514]*kernel[7]+tmp[1515]*kernel[8];
				ans[1415]<=tmp[1314]*kernel[0]+tmp[1315]*kernel[1]+tmp[1316]*kernel[2]+tmp[1414]*kernel[3]+tmp[1415]*kernel[4]+tmp[1416]*kernel[5]+tmp[1514]*kernel[6]+tmp[1515]*kernel[7]+tmp[1516]*kernel[8];
				ans[1416]<=tmp[1315]*kernel[0]+tmp[1316]*kernel[1]+tmp[1317]*kernel[2]+tmp[1415]*kernel[3]+tmp[1416]*kernel[4]+tmp[1417]*kernel[5]+tmp[1515]*kernel[6]+tmp[1516]*kernel[7]+tmp[1517]*kernel[8];
				ans[1417]<=tmp[1316]*kernel[0]+tmp[1317]*kernel[1]+tmp[1318]*kernel[2]+tmp[1416]*kernel[3]+tmp[1417]*kernel[4]+tmp[1418]*kernel[5]+tmp[1516]*kernel[6]+tmp[1517]*kernel[7]+tmp[1518]*kernel[8];
				ans[1418]<=tmp[1317]*kernel[0]+tmp[1318]*kernel[1]+tmp[1319]*kernel[2]+tmp[1417]*kernel[3]+tmp[1418]*kernel[4]+tmp[1419]*kernel[5]+tmp[1517]*kernel[6]+tmp[1518]*kernel[7]+tmp[1519]*kernel[8];
				ans[1419]<=tmp[1318]*kernel[0]+tmp[1319]*kernel[1]+tmp[1320]*kernel[2]+tmp[1418]*kernel[3]+tmp[1419]*kernel[4]+tmp[1420]*kernel[5]+tmp[1518]*kernel[6]+tmp[1519]*kernel[7]+tmp[1520]*kernel[8];
				ans[1420]<=tmp[1319]*kernel[0]+tmp[1320]*kernel[1]+tmp[1321]*kernel[2]+tmp[1419]*kernel[3]+tmp[1420]*kernel[4]+tmp[1421]*kernel[5]+tmp[1519]*kernel[6]+tmp[1520]*kernel[7]+tmp[1521]*kernel[8];
				ans[1421]<=tmp[1320]*kernel[0]+tmp[1321]*kernel[1]+tmp[1322]*kernel[2]+tmp[1420]*kernel[3]+tmp[1421]*kernel[4]+tmp[1422]*kernel[5]+tmp[1520]*kernel[6]+tmp[1521]*kernel[7]+tmp[1522]*kernel[8];
				ans[1422]<=tmp[1321]*kernel[0]+tmp[1322]*kernel[1]+tmp[1323]*kernel[2]+tmp[1421]*kernel[3]+tmp[1422]*kernel[4]+tmp[1423]*kernel[5]+tmp[1521]*kernel[6]+tmp[1522]*kernel[7]+tmp[1523]*kernel[8];
				ans[1423]<=tmp[1322]*kernel[0]+tmp[1323]*kernel[1]+tmp[1324]*kernel[2]+tmp[1422]*kernel[3]+tmp[1423]*kernel[4]+tmp[1424]*kernel[5]+tmp[1522]*kernel[6]+tmp[1523]*kernel[7]+tmp[1524]*kernel[8];
				ans[1424]<=tmp[1323]*kernel[0]+tmp[1324]*kernel[1]+tmp[1325]*kernel[2]+tmp[1423]*kernel[3]+tmp[1424]*kernel[4]+tmp[1425]*kernel[5]+tmp[1523]*kernel[6]+tmp[1524]*kernel[7]+tmp[1525]*kernel[8];
				ans[1425]<=tmp[1324]*kernel[0]+tmp[1325]*kernel[1]+tmp[1326]*kernel[2]+tmp[1424]*kernel[3]+tmp[1425]*kernel[4]+tmp[1426]*kernel[5]+tmp[1524]*kernel[6]+tmp[1525]*kernel[7]+tmp[1526]*kernel[8];
				ans[1426]<=tmp[1325]*kernel[0]+tmp[1326]*kernel[1]+tmp[1327]*kernel[2]+tmp[1425]*kernel[3]+tmp[1426]*kernel[4]+tmp[1427]*kernel[5]+tmp[1525]*kernel[6]+tmp[1526]*kernel[7]+tmp[1527]*kernel[8];
				ans[1427]<=tmp[1326]*kernel[0]+tmp[1327]*kernel[1]+tmp[1328]*kernel[2]+tmp[1426]*kernel[3]+tmp[1427]*kernel[4]+tmp[1428]*kernel[5]+tmp[1526]*kernel[6]+tmp[1527]*kernel[7]+tmp[1528]*kernel[8];
				ans[1428]<=tmp[1327]*kernel[0]+tmp[1328]*kernel[1]+tmp[1329]*kernel[2]+tmp[1427]*kernel[3]+tmp[1428]*kernel[4]+tmp[1429]*kernel[5]+tmp[1527]*kernel[6]+tmp[1528]*kernel[7]+tmp[1529]*kernel[8];
				ans[1429]<=tmp[1328]*kernel[0]+tmp[1329]*kernel[1]+tmp[1330]*kernel[2]+tmp[1428]*kernel[3]+tmp[1429]*kernel[4]+tmp[1430]*kernel[5]+tmp[1528]*kernel[6]+tmp[1529]*kernel[7]+tmp[1530]*kernel[8];
				ans[1430]<=tmp[1329]*kernel[0]+tmp[1330]*kernel[1]+tmp[1331]*kernel[2]+tmp[1429]*kernel[3]+tmp[1430]*kernel[4]+tmp[1431]*kernel[5]+tmp[1529]*kernel[6]+tmp[1530]*kernel[7]+tmp[1531]*kernel[8];
				ans[1431]<=tmp[1330]*kernel[0]+tmp[1331]*kernel[1]+tmp[1332]*kernel[2]+tmp[1430]*kernel[3]+tmp[1431]*kernel[4]+tmp[1432]*kernel[5]+tmp[1530]*kernel[6]+tmp[1531]*kernel[7]+tmp[1532]*kernel[8];
				ans[1432]<=tmp[1331]*kernel[0]+tmp[1332]*kernel[1]+tmp[1333]*kernel[2]+tmp[1431]*kernel[3]+tmp[1432]*kernel[4]+tmp[1433]*kernel[5]+tmp[1531]*kernel[6]+tmp[1532]*kernel[7]+tmp[1533]*kernel[8];
				ans[1433]<=tmp[1332]*kernel[0]+tmp[1333]*kernel[1]+tmp[1334]*kernel[2]+tmp[1432]*kernel[3]+tmp[1433]*kernel[4]+tmp[1434]*kernel[5]+tmp[1532]*kernel[6]+tmp[1533]*kernel[7]+tmp[1534]*kernel[8];
				ans[1434]<=tmp[1333]*kernel[0]+tmp[1334]*kernel[1]+tmp[1335]*kernel[2]+tmp[1433]*kernel[3]+tmp[1434]*kernel[4]+tmp[1435]*kernel[5]+tmp[1533]*kernel[6]+tmp[1534]*kernel[7]+tmp[1535]*kernel[8];
				ans[1435]<=tmp[1334]*kernel[0]+tmp[1335]*kernel[1]+tmp[1336]*kernel[2]+tmp[1434]*kernel[3]+tmp[1435]*kernel[4]+tmp[1436]*kernel[5]+tmp[1534]*kernel[6]+tmp[1535]*kernel[7]+tmp[1536]*kernel[8];
				ans[1436]<=tmp[1335]*kernel[0]+tmp[1336]*kernel[1]+tmp[1337]*kernel[2]+tmp[1435]*kernel[3]+tmp[1436]*kernel[4]+tmp[1437]*kernel[5]+tmp[1535]*kernel[6]+tmp[1536]*kernel[7]+tmp[1537]*kernel[8];
				ans[1437]<=tmp[1336]*kernel[0]+tmp[1337]*kernel[1]+tmp[1338]*kernel[2]+tmp[1436]*kernel[3]+tmp[1437]*kernel[4]+tmp[1438]*kernel[5]+tmp[1536]*kernel[6]+tmp[1537]*kernel[7]+tmp[1538]*kernel[8];
				ans[1438]<=tmp[1337]*kernel[0]+tmp[1338]*kernel[1]+tmp[1339]*kernel[2]+tmp[1437]*kernel[3]+tmp[1438]*kernel[4]+tmp[1439]*kernel[5]+tmp[1537]*kernel[6]+tmp[1538]*kernel[7]+tmp[1539]*kernel[8];
				ans[1439]<=tmp[1338]*kernel[0]+tmp[1339]*kernel[1]+tmp[1340]*kernel[2]+tmp[1438]*kernel[3]+tmp[1439]*kernel[4]+tmp[1440]*kernel[5]+tmp[1538]*kernel[6]+tmp[1539]*kernel[7]+tmp[1540]*kernel[8];
				ans[1440]<=tmp[1339]*kernel[0]+tmp[1340]*kernel[1]+tmp[1341]*kernel[2]+tmp[1439]*kernel[3]+tmp[1440]*kernel[4]+tmp[1441]*kernel[5]+tmp[1539]*kernel[6]+tmp[1540]*kernel[7]+tmp[1541]*kernel[8];
				ans[1441]<=tmp[1340]*kernel[0]+tmp[1341]*kernel[1]+tmp[1342]*kernel[2]+tmp[1440]*kernel[3]+tmp[1441]*kernel[4]+tmp[1442]*kernel[5]+tmp[1540]*kernel[6]+tmp[1541]*kernel[7]+tmp[1542]*kernel[8];
				ans[1442]<=tmp[1341]*kernel[0]+tmp[1342]*kernel[1]+tmp[1343]*kernel[2]+tmp[1441]*kernel[3]+tmp[1442]*kernel[4]+tmp[1443]*kernel[5]+tmp[1541]*kernel[6]+tmp[1542]*kernel[7]+tmp[1543]*kernel[8];
				ans[1443]<=tmp[1342]*kernel[0]+tmp[1343]*kernel[1]+tmp[1344]*kernel[2]+tmp[1442]*kernel[3]+tmp[1443]*kernel[4]+tmp[1444]*kernel[5]+tmp[1542]*kernel[6]+tmp[1543]*kernel[7]+tmp[1544]*kernel[8];
				ans[1444]<=tmp[1343]*kernel[0]+tmp[1344]*kernel[1]+tmp[1345]*kernel[2]+tmp[1443]*kernel[3]+tmp[1444]*kernel[4]+tmp[1445]*kernel[5]+tmp[1543]*kernel[6]+tmp[1544]*kernel[7]+tmp[1545]*kernel[8];
				ans[1445]<=tmp[1344]*kernel[0]+tmp[1345]*kernel[1]+tmp[1346]*kernel[2]+tmp[1444]*kernel[3]+tmp[1445]*kernel[4]+tmp[1446]*kernel[5]+tmp[1544]*kernel[6]+tmp[1545]*kernel[7]+tmp[1546]*kernel[8];
				ans[1446]<=tmp[1345]*kernel[0]+tmp[1346]*kernel[1]+tmp[1347]*kernel[2]+tmp[1445]*kernel[3]+tmp[1446]*kernel[4]+tmp[1447]*kernel[5]+tmp[1545]*kernel[6]+tmp[1546]*kernel[7]+tmp[1547]*kernel[8];
				ans[1447]<=tmp[1346]*kernel[0]+tmp[1347]*kernel[1]+tmp[1348]*kernel[2]+tmp[1446]*kernel[3]+tmp[1447]*kernel[4]+tmp[1448]*kernel[5]+tmp[1546]*kernel[6]+tmp[1547]*kernel[7]+tmp[1548]*kernel[8];
				ans[1448]<=tmp[1347]*kernel[0]+tmp[1348]*kernel[1]+tmp[1349]*kernel[2]+tmp[1447]*kernel[3]+tmp[1448]*kernel[4]+tmp[1449]*kernel[5]+tmp[1547]*kernel[6]+tmp[1548]*kernel[7]+tmp[1549]*kernel[8];
				ans[1449]<=tmp[1348]*kernel[0]+tmp[1349]*kernel[1]+tmp[1350]*kernel[2]+tmp[1448]*kernel[3]+tmp[1449]*kernel[4]+tmp[1450]*kernel[5]+tmp[1548]*kernel[6]+tmp[1549]*kernel[7]+tmp[1550]*kernel[8];
				ans[1450]<=tmp[1349]*kernel[0]+tmp[1350]*kernel[1]+tmp[1351]*kernel[2]+tmp[1449]*kernel[3]+tmp[1450]*kernel[4]+tmp[1451]*kernel[5]+tmp[1549]*kernel[6]+tmp[1550]*kernel[7]+tmp[1551]*kernel[8];
				ans[1451]<=tmp[1350]*kernel[0]+tmp[1351]*kernel[1]+tmp[1352]*kernel[2]+tmp[1450]*kernel[3]+tmp[1451]*kernel[4]+tmp[1452]*kernel[5]+tmp[1550]*kernel[6]+tmp[1551]*kernel[7]+tmp[1552]*kernel[8];
				ans[1452]<=tmp[1351]*kernel[0]+tmp[1352]*kernel[1]+tmp[1353]*kernel[2]+tmp[1451]*kernel[3]+tmp[1452]*kernel[4]+tmp[1453]*kernel[5]+tmp[1551]*kernel[6]+tmp[1552]*kernel[7]+tmp[1553]*kernel[8];
				ans[1453]<=tmp[1352]*kernel[0]+tmp[1353]*kernel[1]+tmp[1354]*kernel[2]+tmp[1452]*kernel[3]+tmp[1453]*kernel[4]+tmp[1454]*kernel[5]+tmp[1552]*kernel[6]+tmp[1553]*kernel[7]+tmp[1554]*kernel[8];
				ans[1454]<=tmp[1353]*kernel[0]+tmp[1354]*kernel[1]+tmp[1355]*kernel[2]+tmp[1453]*kernel[3]+tmp[1454]*kernel[4]+tmp[1455]*kernel[5]+tmp[1553]*kernel[6]+tmp[1554]*kernel[7]+tmp[1555]*kernel[8];
				ans[1455]<=tmp[1354]*kernel[0]+tmp[1355]*kernel[1]+tmp[1356]*kernel[2]+tmp[1454]*kernel[3]+tmp[1455]*kernel[4]+tmp[1456]*kernel[5]+tmp[1554]*kernel[6]+tmp[1555]*kernel[7]+tmp[1556]*kernel[8];
				ans[1456]<=tmp[1355]*kernel[0]+tmp[1356]*kernel[1]+tmp[1357]*kernel[2]+tmp[1455]*kernel[3]+tmp[1456]*kernel[4]+tmp[1457]*kernel[5]+tmp[1555]*kernel[6]+tmp[1556]*kernel[7]+tmp[1557]*kernel[8];
				ans[1457]<=tmp[1356]*kernel[0]+tmp[1357]*kernel[1]+tmp[1358]*kernel[2]+tmp[1456]*kernel[3]+tmp[1457]*kernel[4]+tmp[1458]*kernel[5]+tmp[1556]*kernel[6]+tmp[1557]*kernel[7]+tmp[1558]*kernel[8];
				ans[1458]<=tmp[1357]*kernel[0]+tmp[1358]*kernel[1]+tmp[1359]*kernel[2]+tmp[1457]*kernel[3]+tmp[1458]*kernel[4]+tmp[1459]*kernel[5]+tmp[1557]*kernel[6]+tmp[1558]*kernel[7]+tmp[1559]*kernel[8];
				ans[1459]<=tmp[1358]*kernel[0]+tmp[1359]*kernel[1]+tmp[1360]*kernel[2]+tmp[1458]*kernel[3]+tmp[1459]*kernel[4]+tmp[1460]*kernel[5]+tmp[1558]*kernel[6]+tmp[1559]*kernel[7]+tmp[1560]*kernel[8];
				ans[1460]<=tmp[1359]*kernel[0]+tmp[1360]*kernel[1]+tmp[1361]*kernel[2]+tmp[1459]*kernel[3]+tmp[1460]*kernel[4]+tmp[1461]*kernel[5]+tmp[1559]*kernel[6]+tmp[1560]*kernel[7]+tmp[1561]*kernel[8];
				ans[1461]<=tmp[1360]*kernel[0]+tmp[1361]*kernel[1]+tmp[1362]*kernel[2]+tmp[1460]*kernel[3]+tmp[1461]*kernel[4]+tmp[1462]*kernel[5]+tmp[1560]*kernel[6]+tmp[1561]*kernel[7]+tmp[1562]*kernel[8];
				ans[1462]<=tmp[1361]*kernel[0]+tmp[1362]*kernel[1]+tmp[1363]*kernel[2]+tmp[1461]*kernel[3]+tmp[1462]*kernel[4]+tmp[1463]*kernel[5]+tmp[1561]*kernel[6]+tmp[1562]*kernel[7]+tmp[1563]*kernel[8];
				ans[1463]<=tmp[1362]*kernel[0]+tmp[1363]*kernel[1]+tmp[1364]*kernel[2]+tmp[1462]*kernel[3]+tmp[1463]*kernel[4]+tmp[1464]*kernel[5]+tmp[1562]*kernel[6]+tmp[1563]*kernel[7]+tmp[1564]*kernel[8];
				ans[1464]<=tmp[1363]*kernel[0]+tmp[1364]*kernel[1]+tmp[1365]*kernel[2]+tmp[1463]*kernel[3]+tmp[1464]*kernel[4]+tmp[1465]*kernel[5]+tmp[1563]*kernel[6]+tmp[1564]*kernel[7]+tmp[1565]*kernel[8];
				ans[1465]<=tmp[1364]*kernel[0]+tmp[1365]*kernel[1]+tmp[1366]*kernel[2]+tmp[1464]*kernel[3]+tmp[1465]*kernel[4]+tmp[1466]*kernel[5]+tmp[1564]*kernel[6]+tmp[1565]*kernel[7]+tmp[1566]*kernel[8];
				ans[1466]<=tmp[1365]*kernel[0]+tmp[1366]*kernel[1]+tmp[1367]*kernel[2]+tmp[1465]*kernel[3]+tmp[1466]*kernel[4]+tmp[1467]*kernel[5]+tmp[1565]*kernel[6]+tmp[1566]*kernel[7]+tmp[1567]*kernel[8];
				ans[1467]<=tmp[1366]*kernel[0]+tmp[1367]*kernel[1]+tmp[1368]*kernel[2]+tmp[1466]*kernel[3]+tmp[1467]*kernel[4]+tmp[1468]*kernel[5]+tmp[1566]*kernel[6]+tmp[1567]*kernel[7]+tmp[1568]*kernel[8];
				ans[1468]<=tmp[1367]*kernel[0]+tmp[1368]*kernel[1]+tmp[1369]*kernel[2]+tmp[1467]*kernel[3]+tmp[1468]*kernel[4]+tmp[1469]*kernel[5]+tmp[1567]*kernel[6]+tmp[1568]*kernel[7]+tmp[1569]*kernel[8];
				ans[1469]<=tmp[1368]*kernel[0]+tmp[1369]*kernel[1]+tmp[1370]*kernel[2]+tmp[1468]*kernel[3]+tmp[1469]*kernel[4]+tmp[1470]*kernel[5]+tmp[1568]*kernel[6]+tmp[1569]*kernel[7]+tmp[1570]*kernel[8];
				ans[1470]<=tmp[1369]*kernel[0]+tmp[1370]*kernel[1]+tmp[1371]*kernel[2]+tmp[1469]*kernel[3]+tmp[1470]*kernel[4]+tmp[1471]*kernel[5]+tmp[1569]*kernel[6]+tmp[1570]*kernel[7]+tmp[1571]*kernel[8];
				ans[1471]<=tmp[1370]*kernel[0]+tmp[1371]*kernel[1]+tmp[1372]*kernel[2]+tmp[1470]*kernel[3]+tmp[1471]*kernel[4]+tmp[1472]*kernel[5]+tmp[1570]*kernel[6]+tmp[1571]*kernel[7]+tmp[1572]*kernel[8];
				ans[1472]<=tmp[1371]*kernel[0]+tmp[1372]*kernel[1]+tmp[1373]*kernel[2]+tmp[1471]*kernel[3]+tmp[1472]*kernel[4]+tmp[1473]*kernel[5]+tmp[1571]*kernel[6]+tmp[1572]*kernel[7]+tmp[1573]*kernel[8];
				ans[1473]<=tmp[1372]*kernel[0]+tmp[1373]*kernel[1]+tmp[1374]*kernel[2]+tmp[1472]*kernel[3]+tmp[1473]*kernel[4]+tmp[1474]*kernel[5]+tmp[1572]*kernel[6]+tmp[1573]*kernel[7]+tmp[1574]*kernel[8];
				ans[1474]<=tmp[1373]*kernel[0]+tmp[1374]*kernel[1]+tmp[1375]*kernel[2]+tmp[1473]*kernel[3]+tmp[1474]*kernel[4]+tmp[1475]*kernel[5]+tmp[1573]*kernel[6]+tmp[1574]*kernel[7]+tmp[1575]*kernel[8];
				ans[1475]<=tmp[1374]*kernel[0]+tmp[1375]*kernel[1]+tmp[1376]*kernel[2]+tmp[1474]*kernel[3]+tmp[1475]*kernel[4]+tmp[1476]*kernel[5]+tmp[1574]*kernel[6]+tmp[1575]*kernel[7]+tmp[1576]*kernel[8];
				ans[1476]<=tmp[1375]*kernel[0]+tmp[1376]*kernel[1]+tmp[1377]*kernel[2]+tmp[1475]*kernel[3]+tmp[1476]*kernel[4]+tmp[1477]*kernel[5]+tmp[1575]*kernel[6]+tmp[1576]*kernel[7]+tmp[1577]*kernel[8];
				ans[1477]<=tmp[1376]*kernel[0]+tmp[1377]*kernel[1]+tmp[1378]*kernel[2]+tmp[1476]*kernel[3]+tmp[1477]*kernel[4]+tmp[1478]*kernel[5]+tmp[1576]*kernel[6]+tmp[1577]*kernel[7]+tmp[1578]*kernel[8];
				ans[1478]<=tmp[1377]*kernel[0]+tmp[1378]*kernel[1]+tmp[1379]*kernel[2]+tmp[1477]*kernel[3]+tmp[1478]*kernel[4]+tmp[1479]*kernel[5]+tmp[1577]*kernel[6]+tmp[1578]*kernel[7]+tmp[1579]*kernel[8];
				ans[1479]<=tmp[1378]*kernel[0]+tmp[1379]*kernel[1]+tmp[1380]*kernel[2]+tmp[1478]*kernel[3]+tmp[1479]*kernel[4]+tmp[1480]*kernel[5]+tmp[1578]*kernel[6]+tmp[1579]*kernel[7]+tmp[1580]*kernel[8];
				ans[1480]<=tmp[1379]*kernel[0]+tmp[1380]*kernel[1]+tmp[1381]*kernel[2]+tmp[1479]*kernel[3]+tmp[1480]*kernel[4]+tmp[1481]*kernel[5]+tmp[1579]*kernel[6]+tmp[1580]*kernel[7]+tmp[1581]*kernel[8];
				ans[1481]<=tmp[1380]*kernel[0]+tmp[1381]*kernel[1]+tmp[1382]*kernel[2]+tmp[1480]*kernel[3]+tmp[1481]*kernel[4]+tmp[1482]*kernel[5]+tmp[1580]*kernel[6]+tmp[1581]*kernel[7]+tmp[1582]*kernel[8];
				ans[1482]<=tmp[1381]*kernel[0]+tmp[1382]*kernel[1]+tmp[1383]*kernel[2]+tmp[1481]*kernel[3]+tmp[1482]*kernel[4]+tmp[1483]*kernel[5]+tmp[1581]*kernel[6]+tmp[1582]*kernel[7]+tmp[1583]*kernel[8];
				ans[1483]<=tmp[1382]*kernel[0]+tmp[1383]*kernel[1]+tmp[1384]*kernel[2]+tmp[1482]*kernel[3]+tmp[1483]*kernel[4]+tmp[1484]*kernel[5]+tmp[1582]*kernel[6]+tmp[1583]*kernel[7]+tmp[1584]*kernel[8];
				ans[1484]<=tmp[1383]*kernel[0]+tmp[1384]*kernel[1]+tmp[1385]*kernel[2]+tmp[1483]*kernel[3]+tmp[1484]*kernel[4]+tmp[1485]*kernel[5]+tmp[1583]*kernel[6]+tmp[1584]*kernel[7]+tmp[1585]*kernel[8];
				ans[1485]<=tmp[1384]*kernel[0]+tmp[1385]*kernel[1]+tmp[1386]*kernel[2]+tmp[1484]*kernel[3]+tmp[1485]*kernel[4]+tmp[1486]*kernel[5]+tmp[1584]*kernel[6]+tmp[1585]*kernel[7]+tmp[1586]*kernel[8];
				ans[1486]<=tmp[1385]*kernel[0]+tmp[1386]*kernel[1]+tmp[1387]*kernel[2]+tmp[1485]*kernel[3]+tmp[1486]*kernel[4]+tmp[1487]*kernel[5]+tmp[1585]*kernel[6]+tmp[1586]*kernel[7]+tmp[1587]*kernel[8];
				ans[1487]<=tmp[1386]*kernel[0]+tmp[1387]*kernel[1]+tmp[1388]*kernel[2]+tmp[1486]*kernel[3]+tmp[1487]*kernel[4]+tmp[1488]*kernel[5]+tmp[1586]*kernel[6]+tmp[1587]*kernel[7]+tmp[1588]*kernel[8];
				ans[1488]<=tmp[1387]*kernel[0]+tmp[1388]*kernel[1]+tmp[1389]*kernel[2]+tmp[1487]*kernel[3]+tmp[1488]*kernel[4]+tmp[1489]*kernel[5]+tmp[1587]*kernel[6]+tmp[1588]*kernel[7]+tmp[1589]*kernel[8];
				ans[1489]<=tmp[1388]*kernel[0]+tmp[1389]*kernel[1]+tmp[1390]*kernel[2]+tmp[1488]*kernel[3]+tmp[1489]*kernel[4]+tmp[1490]*kernel[5]+tmp[1588]*kernel[6]+tmp[1589]*kernel[7]+tmp[1590]*kernel[8];
				ans[1490]<=tmp[1389]*kernel[0]+tmp[1390]*kernel[1]+tmp[1391]*kernel[2]+tmp[1489]*kernel[3]+tmp[1490]*kernel[4]+tmp[1491]*kernel[5]+tmp[1589]*kernel[6]+tmp[1590]*kernel[7]+tmp[1591]*kernel[8];
				ans[1491]<=tmp[1390]*kernel[0]+tmp[1391]*kernel[1]+tmp[1392]*kernel[2]+tmp[1490]*kernel[3]+tmp[1491]*kernel[4]+tmp[1492]*kernel[5]+tmp[1590]*kernel[6]+tmp[1591]*kernel[7]+tmp[1592]*kernel[8];
				ans[1492]<=tmp[1391]*kernel[0]+tmp[1392]*kernel[1]+tmp[1393]*kernel[2]+tmp[1491]*kernel[3]+tmp[1492]*kernel[4]+tmp[1493]*kernel[5]+tmp[1591]*kernel[6]+tmp[1592]*kernel[7]+tmp[1593]*kernel[8];
				ans[1493]<=tmp[1392]*kernel[0]+tmp[1393]*kernel[1]+tmp[1394]*kernel[2]+tmp[1492]*kernel[3]+tmp[1493]*kernel[4]+tmp[1494]*kernel[5]+tmp[1592]*kernel[6]+tmp[1593]*kernel[7]+tmp[1594]*kernel[8];
				ans[1494]<=tmp[1393]*kernel[0]+tmp[1394]*kernel[1]+tmp[1395]*kernel[2]+tmp[1493]*kernel[3]+tmp[1494]*kernel[4]+tmp[1495]*kernel[5]+tmp[1593]*kernel[6]+tmp[1594]*kernel[7]+tmp[1595]*kernel[8];
				ans[1495]<=tmp[1394]*kernel[0]+tmp[1395]*kernel[1]+tmp[1396]*kernel[2]+tmp[1494]*kernel[3]+tmp[1495]*kernel[4]+tmp[1496]*kernel[5]+tmp[1594]*kernel[6]+tmp[1595]*kernel[7]+tmp[1596]*kernel[8];
				ans[1496]<=tmp[1395]*kernel[0]+tmp[1396]*kernel[1]+tmp[1397]*kernel[2]+tmp[1495]*kernel[3]+tmp[1496]*kernel[4]+tmp[1497]*kernel[5]+tmp[1595]*kernel[6]+tmp[1596]*kernel[7]+tmp[1597]*kernel[8];
				ans[1497]<=tmp[1396]*kernel[0]+tmp[1397]*kernel[1]+tmp[1398]*kernel[2]+tmp[1496]*kernel[3]+tmp[1497]*kernel[4]+tmp[1498]*kernel[5]+tmp[1596]*kernel[6]+tmp[1597]*kernel[7]+tmp[1598]*kernel[8];
				ans[1498]<=tmp[1397]*kernel[0]+tmp[1398]*kernel[1]+tmp[1399]*kernel[2]+tmp[1497]*kernel[3]+tmp[1498]*kernel[4]+tmp[1499]*kernel[5]+tmp[1597]*kernel[6]+tmp[1598]*kernel[7]+tmp[1599]*kernel[8];
				ans[1499]<=tmp[1398]*kernel[0]+tmp[1399]*kernel[1]+tmp[1498]*kernel[3]+tmp[1499]*kernel[4]+tmp[1598]*kernel[6]+tmp[1599]*kernel[7];
				ans[1500]<=tmp[1400]*kernel[1]+tmp[1401]*kernel[2]+tmp[1500]*kernel[4]+tmp[1501]*kernel[5]+tmp[1600]*kernel[7]+tmp[1601]*kernel[8];
				ans[1501]<=tmp[1400]*kernel[0]+tmp[1401]*kernel[1]+tmp[1402]*kernel[2]+tmp[1500]*kernel[3]+tmp[1501]*kernel[4]+tmp[1502]*kernel[5]+tmp[1600]*kernel[6]+tmp[1601]*kernel[7]+tmp[1602]*kernel[8];
				ans[1502]<=tmp[1401]*kernel[0]+tmp[1402]*kernel[1]+tmp[1403]*kernel[2]+tmp[1501]*kernel[3]+tmp[1502]*kernel[4]+tmp[1503]*kernel[5]+tmp[1601]*kernel[6]+tmp[1602]*kernel[7]+tmp[1603]*kernel[8];
				ans[1503]<=tmp[1402]*kernel[0]+tmp[1403]*kernel[1]+tmp[1404]*kernel[2]+tmp[1502]*kernel[3]+tmp[1503]*kernel[4]+tmp[1504]*kernel[5]+tmp[1602]*kernel[6]+tmp[1603]*kernel[7]+tmp[1604]*kernel[8];
				ans[1504]<=tmp[1403]*kernel[0]+tmp[1404]*kernel[1]+tmp[1405]*kernel[2]+tmp[1503]*kernel[3]+tmp[1504]*kernel[4]+tmp[1505]*kernel[5]+tmp[1603]*kernel[6]+tmp[1604]*kernel[7]+tmp[1605]*kernel[8];
				ans[1505]<=tmp[1404]*kernel[0]+tmp[1405]*kernel[1]+tmp[1406]*kernel[2]+tmp[1504]*kernel[3]+tmp[1505]*kernel[4]+tmp[1506]*kernel[5]+tmp[1604]*kernel[6]+tmp[1605]*kernel[7]+tmp[1606]*kernel[8];
				ans[1506]<=tmp[1405]*kernel[0]+tmp[1406]*kernel[1]+tmp[1407]*kernel[2]+tmp[1505]*kernel[3]+tmp[1506]*kernel[4]+tmp[1507]*kernel[5]+tmp[1605]*kernel[6]+tmp[1606]*kernel[7]+tmp[1607]*kernel[8];
				ans[1507]<=tmp[1406]*kernel[0]+tmp[1407]*kernel[1]+tmp[1408]*kernel[2]+tmp[1506]*kernel[3]+tmp[1507]*kernel[4]+tmp[1508]*kernel[5]+tmp[1606]*kernel[6]+tmp[1607]*kernel[7]+tmp[1608]*kernel[8];
				ans[1508]<=tmp[1407]*kernel[0]+tmp[1408]*kernel[1]+tmp[1409]*kernel[2]+tmp[1507]*kernel[3]+tmp[1508]*kernel[4]+tmp[1509]*kernel[5]+tmp[1607]*kernel[6]+tmp[1608]*kernel[7]+tmp[1609]*kernel[8];
				ans[1509]<=tmp[1408]*kernel[0]+tmp[1409]*kernel[1]+tmp[1410]*kernel[2]+tmp[1508]*kernel[3]+tmp[1509]*kernel[4]+tmp[1510]*kernel[5]+tmp[1608]*kernel[6]+tmp[1609]*kernel[7]+tmp[1610]*kernel[8];
				ans[1510]<=tmp[1409]*kernel[0]+tmp[1410]*kernel[1]+tmp[1411]*kernel[2]+tmp[1509]*kernel[3]+tmp[1510]*kernel[4]+tmp[1511]*kernel[5]+tmp[1609]*kernel[6]+tmp[1610]*kernel[7]+tmp[1611]*kernel[8];
				ans[1511]<=tmp[1410]*kernel[0]+tmp[1411]*kernel[1]+tmp[1412]*kernel[2]+tmp[1510]*kernel[3]+tmp[1511]*kernel[4]+tmp[1512]*kernel[5]+tmp[1610]*kernel[6]+tmp[1611]*kernel[7]+tmp[1612]*kernel[8];
				ans[1512]<=tmp[1411]*kernel[0]+tmp[1412]*kernel[1]+tmp[1413]*kernel[2]+tmp[1511]*kernel[3]+tmp[1512]*kernel[4]+tmp[1513]*kernel[5]+tmp[1611]*kernel[6]+tmp[1612]*kernel[7]+tmp[1613]*kernel[8];
				ans[1513]<=tmp[1412]*kernel[0]+tmp[1413]*kernel[1]+tmp[1414]*kernel[2]+tmp[1512]*kernel[3]+tmp[1513]*kernel[4]+tmp[1514]*kernel[5]+tmp[1612]*kernel[6]+tmp[1613]*kernel[7]+tmp[1614]*kernel[8];
				ans[1514]<=tmp[1413]*kernel[0]+tmp[1414]*kernel[1]+tmp[1415]*kernel[2]+tmp[1513]*kernel[3]+tmp[1514]*kernel[4]+tmp[1515]*kernel[5]+tmp[1613]*kernel[6]+tmp[1614]*kernel[7]+tmp[1615]*kernel[8];
				ans[1515]<=tmp[1414]*kernel[0]+tmp[1415]*kernel[1]+tmp[1416]*kernel[2]+tmp[1514]*kernel[3]+tmp[1515]*kernel[4]+tmp[1516]*kernel[5]+tmp[1614]*kernel[6]+tmp[1615]*kernel[7]+tmp[1616]*kernel[8];
				ans[1516]<=tmp[1415]*kernel[0]+tmp[1416]*kernel[1]+tmp[1417]*kernel[2]+tmp[1515]*kernel[3]+tmp[1516]*kernel[4]+tmp[1517]*kernel[5]+tmp[1615]*kernel[6]+tmp[1616]*kernel[7]+tmp[1617]*kernel[8];
				ans[1517]<=tmp[1416]*kernel[0]+tmp[1417]*kernel[1]+tmp[1418]*kernel[2]+tmp[1516]*kernel[3]+tmp[1517]*kernel[4]+tmp[1518]*kernel[5]+tmp[1616]*kernel[6]+tmp[1617]*kernel[7]+tmp[1618]*kernel[8];
				ans[1518]<=tmp[1417]*kernel[0]+tmp[1418]*kernel[1]+tmp[1419]*kernel[2]+tmp[1517]*kernel[3]+tmp[1518]*kernel[4]+tmp[1519]*kernel[5]+tmp[1617]*kernel[6]+tmp[1618]*kernel[7]+tmp[1619]*kernel[8];
				ans[1519]<=tmp[1418]*kernel[0]+tmp[1419]*kernel[1]+tmp[1420]*kernel[2]+tmp[1518]*kernel[3]+tmp[1519]*kernel[4]+tmp[1520]*kernel[5]+tmp[1618]*kernel[6]+tmp[1619]*kernel[7]+tmp[1620]*kernel[8];
				ans[1520]<=tmp[1419]*kernel[0]+tmp[1420]*kernel[1]+tmp[1421]*kernel[2]+tmp[1519]*kernel[3]+tmp[1520]*kernel[4]+tmp[1521]*kernel[5]+tmp[1619]*kernel[6]+tmp[1620]*kernel[7]+tmp[1621]*kernel[8];
				ans[1521]<=tmp[1420]*kernel[0]+tmp[1421]*kernel[1]+tmp[1422]*kernel[2]+tmp[1520]*kernel[3]+tmp[1521]*kernel[4]+tmp[1522]*kernel[5]+tmp[1620]*kernel[6]+tmp[1621]*kernel[7]+tmp[1622]*kernel[8];
				ans[1522]<=tmp[1421]*kernel[0]+tmp[1422]*kernel[1]+tmp[1423]*kernel[2]+tmp[1521]*kernel[3]+tmp[1522]*kernel[4]+tmp[1523]*kernel[5]+tmp[1621]*kernel[6]+tmp[1622]*kernel[7]+tmp[1623]*kernel[8];
				ans[1523]<=tmp[1422]*kernel[0]+tmp[1423]*kernel[1]+tmp[1424]*kernel[2]+tmp[1522]*kernel[3]+tmp[1523]*kernel[4]+tmp[1524]*kernel[5]+tmp[1622]*kernel[6]+tmp[1623]*kernel[7]+tmp[1624]*kernel[8];
				ans[1524]<=tmp[1423]*kernel[0]+tmp[1424]*kernel[1]+tmp[1425]*kernel[2]+tmp[1523]*kernel[3]+tmp[1524]*kernel[4]+tmp[1525]*kernel[5]+tmp[1623]*kernel[6]+tmp[1624]*kernel[7]+tmp[1625]*kernel[8];
				ans[1525]<=tmp[1424]*kernel[0]+tmp[1425]*kernel[1]+tmp[1426]*kernel[2]+tmp[1524]*kernel[3]+tmp[1525]*kernel[4]+tmp[1526]*kernel[5]+tmp[1624]*kernel[6]+tmp[1625]*kernel[7]+tmp[1626]*kernel[8];
				ans[1526]<=tmp[1425]*kernel[0]+tmp[1426]*kernel[1]+tmp[1427]*kernel[2]+tmp[1525]*kernel[3]+tmp[1526]*kernel[4]+tmp[1527]*kernel[5]+tmp[1625]*kernel[6]+tmp[1626]*kernel[7]+tmp[1627]*kernel[8];
				ans[1527]<=tmp[1426]*kernel[0]+tmp[1427]*kernel[1]+tmp[1428]*kernel[2]+tmp[1526]*kernel[3]+tmp[1527]*kernel[4]+tmp[1528]*kernel[5]+tmp[1626]*kernel[6]+tmp[1627]*kernel[7]+tmp[1628]*kernel[8];
				ans[1528]<=tmp[1427]*kernel[0]+tmp[1428]*kernel[1]+tmp[1429]*kernel[2]+tmp[1527]*kernel[3]+tmp[1528]*kernel[4]+tmp[1529]*kernel[5]+tmp[1627]*kernel[6]+tmp[1628]*kernel[7]+tmp[1629]*kernel[8];
				ans[1529]<=tmp[1428]*kernel[0]+tmp[1429]*kernel[1]+tmp[1430]*kernel[2]+tmp[1528]*kernel[3]+tmp[1529]*kernel[4]+tmp[1530]*kernel[5]+tmp[1628]*kernel[6]+tmp[1629]*kernel[7]+tmp[1630]*kernel[8];
				ans[1530]<=tmp[1429]*kernel[0]+tmp[1430]*kernel[1]+tmp[1431]*kernel[2]+tmp[1529]*kernel[3]+tmp[1530]*kernel[4]+tmp[1531]*kernel[5]+tmp[1629]*kernel[6]+tmp[1630]*kernel[7]+tmp[1631]*kernel[8];
				ans[1531]<=tmp[1430]*kernel[0]+tmp[1431]*kernel[1]+tmp[1432]*kernel[2]+tmp[1530]*kernel[3]+tmp[1531]*kernel[4]+tmp[1532]*kernel[5]+tmp[1630]*kernel[6]+tmp[1631]*kernel[7]+tmp[1632]*kernel[8];
				ans[1532]<=tmp[1431]*kernel[0]+tmp[1432]*kernel[1]+tmp[1433]*kernel[2]+tmp[1531]*kernel[3]+tmp[1532]*kernel[4]+tmp[1533]*kernel[5]+tmp[1631]*kernel[6]+tmp[1632]*kernel[7]+tmp[1633]*kernel[8];
				ans[1533]<=tmp[1432]*kernel[0]+tmp[1433]*kernel[1]+tmp[1434]*kernel[2]+tmp[1532]*kernel[3]+tmp[1533]*kernel[4]+tmp[1534]*kernel[5]+tmp[1632]*kernel[6]+tmp[1633]*kernel[7]+tmp[1634]*kernel[8];
				ans[1534]<=tmp[1433]*kernel[0]+tmp[1434]*kernel[1]+tmp[1435]*kernel[2]+tmp[1533]*kernel[3]+tmp[1534]*kernel[4]+tmp[1535]*kernel[5]+tmp[1633]*kernel[6]+tmp[1634]*kernel[7]+tmp[1635]*kernel[8];
				ans[1535]<=tmp[1434]*kernel[0]+tmp[1435]*kernel[1]+tmp[1436]*kernel[2]+tmp[1534]*kernel[3]+tmp[1535]*kernel[4]+tmp[1536]*kernel[5]+tmp[1634]*kernel[6]+tmp[1635]*kernel[7]+tmp[1636]*kernel[8];
				ans[1536]<=tmp[1435]*kernel[0]+tmp[1436]*kernel[1]+tmp[1437]*kernel[2]+tmp[1535]*kernel[3]+tmp[1536]*kernel[4]+tmp[1537]*kernel[5]+tmp[1635]*kernel[6]+tmp[1636]*kernel[7]+tmp[1637]*kernel[8];
				ans[1537]<=tmp[1436]*kernel[0]+tmp[1437]*kernel[1]+tmp[1438]*kernel[2]+tmp[1536]*kernel[3]+tmp[1537]*kernel[4]+tmp[1538]*kernel[5]+tmp[1636]*kernel[6]+tmp[1637]*kernel[7]+tmp[1638]*kernel[8];
				ans[1538]<=tmp[1437]*kernel[0]+tmp[1438]*kernel[1]+tmp[1439]*kernel[2]+tmp[1537]*kernel[3]+tmp[1538]*kernel[4]+tmp[1539]*kernel[5]+tmp[1637]*kernel[6]+tmp[1638]*kernel[7]+tmp[1639]*kernel[8];
				ans[1539]<=tmp[1438]*kernel[0]+tmp[1439]*kernel[1]+tmp[1440]*kernel[2]+tmp[1538]*kernel[3]+tmp[1539]*kernel[4]+tmp[1540]*kernel[5]+tmp[1638]*kernel[6]+tmp[1639]*kernel[7]+tmp[1640]*kernel[8];
				ans[1540]<=tmp[1439]*kernel[0]+tmp[1440]*kernel[1]+tmp[1441]*kernel[2]+tmp[1539]*kernel[3]+tmp[1540]*kernel[4]+tmp[1541]*kernel[5]+tmp[1639]*kernel[6]+tmp[1640]*kernel[7]+tmp[1641]*kernel[8];
				ans[1541]<=tmp[1440]*kernel[0]+tmp[1441]*kernel[1]+tmp[1442]*kernel[2]+tmp[1540]*kernel[3]+tmp[1541]*kernel[4]+tmp[1542]*kernel[5]+tmp[1640]*kernel[6]+tmp[1641]*kernel[7]+tmp[1642]*kernel[8];
				ans[1542]<=tmp[1441]*kernel[0]+tmp[1442]*kernel[1]+tmp[1443]*kernel[2]+tmp[1541]*kernel[3]+tmp[1542]*kernel[4]+tmp[1543]*kernel[5]+tmp[1641]*kernel[6]+tmp[1642]*kernel[7]+tmp[1643]*kernel[8];
				ans[1543]<=tmp[1442]*kernel[0]+tmp[1443]*kernel[1]+tmp[1444]*kernel[2]+tmp[1542]*kernel[3]+tmp[1543]*kernel[4]+tmp[1544]*kernel[5]+tmp[1642]*kernel[6]+tmp[1643]*kernel[7]+tmp[1644]*kernel[8];
				ans[1544]<=tmp[1443]*kernel[0]+tmp[1444]*kernel[1]+tmp[1445]*kernel[2]+tmp[1543]*kernel[3]+tmp[1544]*kernel[4]+tmp[1545]*kernel[5]+tmp[1643]*kernel[6]+tmp[1644]*kernel[7]+tmp[1645]*kernel[8];
				ans[1545]<=tmp[1444]*kernel[0]+tmp[1445]*kernel[1]+tmp[1446]*kernel[2]+tmp[1544]*kernel[3]+tmp[1545]*kernel[4]+tmp[1546]*kernel[5]+tmp[1644]*kernel[6]+tmp[1645]*kernel[7]+tmp[1646]*kernel[8];
				ans[1546]<=tmp[1445]*kernel[0]+tmp[1446]*kernel[1]+tmp[1447]*kernel[2]+tmp[1545]*kernel[3]+tmp[1546]*kernel[4]+tmp[1547]*kernel[5]+tmp[1645]*kernel[6]+tmp[1646]*kernel[7]+tmp[1647]*kernel[8];
				ans[1547]<=tmp[1446]*kernel[0]+tmp[1447]*kernel[1]+tmp[1448]*kernel[2]+tmp[1546]*kernel[3]+tmp[1547]*kernel[4]+tmp[1548]*kernel[5]+tmp[1646]*kernel[6]+tmp[1647]*kernel[7]+tmp[1648]*kernel[8];
				ans[1548]<=tmp[1447]*kernel[0]+tmp[1448]*kernel[1]+tmp[1449]*kernel[2]+tmp[1547]*kernel[3]+tmp[1548]*kernel[4]+tmp[1549]*kernel[5]+tmp[1647]*kernel[6]+tmp[1648]*kernel[7]+tmp[1649]*kernel[8];
				ans[1549]<=tmp[1448]*kernel[0]+tmp[1449]*kernel[1]+tmp[1450]*kernel[2]+tmp[1548]*kernel[3]+tmp[1549]*kernel[4]+tmp[1550]*kernel[5]+tmp[1648]*kernel[6]+tmp[1649]*kernel[7]+tmp[1650]*kernel[8];
				ans[1550]<=tmp[1449]*kernel[0]+tmp[1450]*kernel[1]+tmp[1451]*kernel[2]+tmp[1549]*kernel[3]+tmp[1550]*kernel[4]+tmp[1551]*kernel[5]+tmp[1649]*kernel[6]+tmp[1650]*kernel[7]+tmp[1651]*kernel[8];
				ans[1551]<=tmp[1450]*kernel[0]+tmp[1451]*kernel[1]+tmp[1452]*kernel[2]+tmp[1550]*kernel[3]+tmp[1551]*kernel[4]+tmp[1552]*kernel[5]+tmp[1650]*kernel[6]+tmp[1651]*kernel[7]+tmp[1652]*kernel[8];
				ans[1552]<=tmp[1451]*kernel[0]+tmp[1452]*kernel[1]+tmp[1453]*kernel[2]+tmp[1551]*kernel[3]+tmp[1552]*kernel[4]+tmp[1553]*kernel[5]+tmp[1651]*kernel[6]+tmp[1652]*kernel[7]+tmp[1653]*kernel[8];
				ans[1553]<=tmp[1452]*kernel[0]+tmp[1453]*kernel[1]+tmp[1454]*kernel[2]+tmp[1552]*kernel[3]+tmp[1553]*kernel[4]+tmp[1554]*kernel[5]+tmp[1652]*kernel[6]+tmp[1653]*kernel[7]+tmp[1654]*kernel[8];
				ans[1554]<=tmp[1453]*kernel[0]+tmp[1454]*kernel[1]+tmp[1455]*kernel[2]+tmp[1553]*kernel[3]+tmp[1554]*kernel[4]+tmp[1555]*kernel[5]+tmp[1653]*kernel[6]+tmp[1654]*kernel[7]+tmp[1655]*kernel[8];
				ans[1555]<=tmp[1454]*kernel[0]+tmp[1455]*kernel[1]+tmp[1456]*kernel[2]+tmp[1554]*kernel[3]+tmp[1555]*kernel[4]+tmp[1556]*kernel[5]+tmp[1654]*kernel[6]+tmp[1655]*kernel[7]+tmp[1656]*kernel[8];
				ans[1556]<=tmp[1455]*kernel[0]+tmp[1456]*kernel[1]+tmp[1457]*kernel[2]+tmp[1555]*kernel[3]+tmp[1556]*kernel[4]+tmp[1557]*kernel[5]+tmp[1655]*kernel[6]+tmp[1656]*kernel[7]+tmp[1657]*kernel[8];
				ans[1557]<=tmp[1456]*kernel[0]+tmp[1457]*kernel[1]+tmp[1458]*kernel[2]+tmp[1556]*kernel[3]+tmp[1557]*kernel[4]+tmp[1558]*kernel[5]+tmp[1656]*kernel[6]+tmp[1657]*kernel[7]+tmp[1658]*kernel[8];
				ans[1558]<=tmp[1457]*kernel[0]+tmp[1458]*kernel[1]+tmp[1459]*kernel[2]+tmp[1557]*kernel[3]+tmp[1558]*kernel[4]+tmp[1559]*kernel[5]+tmp[1657]*kernel[6]+tmp[1658]*kernel[7]+tmp[1659]*kernel[8];
				ans[1559]<=tmp[1458]*kernel[0]+tmp[1459]*kernel[1]+tmp[1460]*kernel[2]+tmp[1558]*kernel[3]+tmp[1559]*kernel[4]+tmp[1560]*kernel[5]+tmp[1658]*kernel[6]+tmp[1659]*kernel[7]+tmp[1660]*kernel[8];
				ans[1560]<=tmp[1459]*kernel[0]+tmp[1460]*kernel[1]+tmp[1461]*kernel[2]+tmp[1559]*kernel[3]+tmp[1560]*kernel[4]+tmp[1561]*kernel[5]+tmp[1659]*kernel[6]+tmp[1660]*kernel[7]+tmp[1661]*kernel[8];
				ans[1561]<=tmp[1460]*kernel[0]+tmp[1461]*kernel[1]+tmp[1462]*kernel[2]+tmp[1560]*kernel[3]+tmp[1561]*kernel[4]+tmp[1562]*kernel[5]+tmp[1660]*kernel[6]+tmp[1661]*kernel[7]+tmp[1662]*kernel[8];
				ans[1562]<=tmp[1461]*kernel[0]+tmp[1462]*kernel[1]+tmp[1463]*kernel[2]+tmp[1561]*kernel[3]+tmp[1562]*kernel[4]+tmp[1563]*kernel[5]+tmp[1661]*kernel[6]+tmp[1662]*kernel[7]+tmp[1663]*kernel[8];
				ans[1563]<=tmp[1462]*kernel[0]+tmp[1463]*kernel[1]+tmp[1464]*kernel[2]+tmp[1562]*kernel[3]+tmp[1563]*kernel[4]+tmp[1564]*kernel[5]+tmp[1662]*kernel[6]+tmp[1663]*kernel[7]+tmp[1664]*kernel[8];
				ans[1564]<=tmp[1463]*kernel[0]+tmp[1464]*kernel[1]+tmp[1465]*kernel[2]+tmp[1563]*kernel[3]+tmp[1564]*kernel[4]+tmp[1565]*kernel[5]+tmp[1663]*kernel[6]+tmp[1664]*kernel[7]+tmp[1665]*kernel[8];
				ans[1565]<=tmp[1464]*kernel[0]+tmp[1465]*kernel[1]+tmp[1466]*kernel[2]+tmp[1564]*kernel[3]+tmp[1565]*kernel[4]+tmp[1566]*kernel[5]+tmp[1664]*kernel[6]+tmp[1665]*kernel[7]+tmp[1666]*kernel[8];
				ans[1566]<=tmp[1465]*kernel[0]+tmp[1466]*kernel[1]+tmp[1467]*kernel[2]+tmp[1565]*kernel[3]+tmp[1566]*kernel[4]+tmp[1567]*kernel[5]+tmp[1665]*kernel[6]+tmp[1666]*kernel[7]+tmp[1667]*kernel[8];
				ans[1567]<=tmp[1466]*kernel[0]+tmp[1467]*kernel[1]+tmp[1468]*kernel[2]+tmp[1566]*kernel[3]+tmp[1567]*kernel[4]+tmp[1568]*kernel[5]+tmp[1666]*kernel[6]+tmp[1667]*kernel[7]+tmp[1668]*kernel[8];
				ans[1568]<=tmp[1467]*kernel[0]+tmp[1468]*kernel[1]+tmp[1469]*kernel[2]+tmp[1567]*kernel[3]+tmp[1568]*kernel[4]+tmp[1569]*kernel[5]+tmp[1667]*kernel[6]+tmp[1668]*kernel[7]+tmp[1669]*kernel[8];
				ans[1569]<=tmp[1468]*kernel[0]+tmp[1469]*kernel[1]+tmp[1470]*kernel[2]+tmp[1568]*kernel[3]+tmp[1569]*kernel[4]+tmp[1570]*kernel[5]+tmp[1668]*kernel[6]+tmp[1669]*kernel[7]+tmp[1670]*kernel[8];
				ans[1570]<=tmp[1469]*kernel[0]+tmp[1470]*kernel[1]+tmp[1471]*kernel[2]+tmp[1569]*kernel[3]+tmp[1570]*kernel[4]+tmp[1571]*kernel[5]+tmp[1669]*kernel[6]+tmp[1670]*kernel[7]+tmp[1671]*kernel[8];
				ans[1571]<=tmp[1470]*kernel[0]+tmp[1471]*kernel[1]+tmp[1472]*kernel[2]+tmp[1570]*kernel[3]+tmp[1571]*kernel[4]+tmp[1572]*kernel[5]+tmp[1670]*kernel[6]+tmp[1671]*kernel[7]+tmp[1672]*kernel[8];
				ans[1572]<=tmp[1471]*kernel[0]+tmp[1472]*kernel[1]+tmp[1473]*kernel[2]+tmp[1571]*kernel[3]+tmp[1572]*kernel[4]+tmp[1573]*kernel[5]+tmp[1671]*kernel[6]+tmp[1672]*kernel[7]+tmp[1673]*kernel[8];
				ans[1573]<=tmp[1472]*kernel[0]+tmp[1473]*kernel[1]+tmp[1474]*kernel[2]+tmp[1572]*kernel[3]+tmp[1573]*kernel[4]+tmp[1574]*kernel[5]+tmp[1672]*kernel[6]+tmp[1673]*kernel[7]+tmp[1674]*kernel[8];
				ans[1574]<=tmp[1473]*kernel[0]+tmp[1474]*kernel[1]+tmp[1475]*kernel[2]+tmp[1573]*kernel[3]+tmp[1574]*kernel[4]+tmp[1575]*kernel[5]+tmp[1673]*kernel[6]+tmp[1674]*kernel[7]+tmp[1675]*kernel[8];
				ans[1575]<=tmp[1474]*kernel[0]+tmp[1475]*kernel[1]+tmp[1476]*kernel[2]+tmp[1574]*kernel[3]+tmp[1575]*kernel[4]+tmp[1576]*kernel[5]+tmp[1674]*kernel[6]+tmp[1675]*kernel[7]+tmp[1676]*kernel[8];
				ans[1576]<=tmp[1475]*kernel[0]+tmp[1476]*kernel[1]+tmp[1477]*kernel[2]+tmp[1575]*kernel[3]+tmp[1576]*kernel[4]+tmp[1577]*kernel[5]+tmp[1675]*kernel[6]+tmp[1676]*kernel[7]+tmp[1677]*kernel[8];
				ans[1577]<=tmp[1476]*kernel[0]+tmp[1477]*kernel[1]+tmp[1478]*kernel[2]+tmp[1576]*kernel[3]+tmp[1577]*kernel[4]+tmp[1578]*kernel[5]+tmp[1676]*kernel[6]+tmp[1677]*kernel[7]+tmp[1678]*kernel[8];
				ans[1578]<=tmp[1477]*kernel[0]+tmp[1478]*kernel[1]+tmp[1479]*kernel[2]+tmp[1577]*kernel[3]+tmp[1578]*kernel[4]+tmp[1579]*kernel[5]+tmp[1677]*kernel[6]+tmp[1678]*kernel[7]+tmp[1679]*kernel[8];
				ans[1579]<=tmp[1478]*kernel[0]+tmp[1479]*kernel[1]+tmp[1480]*kernel[2]+tmp[1578]*kernel[3]+tmp[1579]*kernel[4]+tmp[1580]*kernel[5]+tmp[1678]*kernel[6]+tmp[1679]*kernel[7]+tmp[1680]*kernel[8];
				ans[1580]<=tmp[1479]*kernel[0]+tmp[1480]*kernel[1]+tmp[1481]*kernel[2]+tmp[1579]*kernel[3]+tmp[1580]*kernel[4]+tmp[1581]*kernel[5]+tmp[1679]*kernel[6]+tmp[1680]*kernel[7]+tmp[1681]*kernel[8];
				ans[1581]<=tmp[1480]*kernel[0]+tmp[1481]*kernel[1]+tmp[1482]*kernel[2]+tmp[1580]*kernel[3]+tmp[1581]*kernel[4]+tmp[1582]*kernel[5]+tmp[1680]*kernel[6]+tmp[1681]*kernel[7]+tmp[1682]*kernel[8];
				ans[1582]<=tmp[1481]*kernel[0]+tmp[1482]*kernel[1]+tmp[1483]*kernel[2]+tmp[1581]*kernel[3]+tmp[1582]*kernel[4]+tmp[1583]*kernel[5]+tmp[1681]*kernel[6]+tmp[1682]*kernel[7]+tmp[1683]*kernel[8];
				ans[1583]<=tmp[1482]*kernel[0]+tmp[1483]*kernel[1]+tmp[1484]*kernel[2]+tmp[1582]*kernel[3]+tmp[1583]*kernel[4]+tmp[1584]*kernel[5]+tmp[1682]*kernel[6]+tmp[1683]*kernel[7]+tmp[1684]*kernel[8];
				ans[1584]<=tmp[1483]*kernel[0]+tmp[1484]*kernel[1]+tmp[1485]*kernel[2]+tmp[1583]*kernel[3]+tmp[1584]*kernel[4]+tmp[1585]*kernel[5]+tmp[1683]*kernel[6]+tmp[1684]*kernel[7]+tmp[1685]*kernel[8];
				ans[1585]<=tmp[1484]*kernel[0]+tmp[1485]*kernel[1]+tmp[1486]*kernel[2]+tmp[1584]*kernel[3]+tmp[1585]*kernel[4]+tmp[1586]*kernel[5]+tmp[1684]*kernel[6]+tmp[1685]*kernel[7]+tmp[1686]*kernel[8];
				ans[1586]<=tmp[1485]*kernel[0]+tmp[1486]*kernel[1]+tmp[1487]*kernel[2]+tmp[1585]*kernel[3]+tmp[1586]*kernel[4]+tmp[1587]*kernel[5]+tmp[1685]*kernel[6]+tmp[1686]*kernel[7]+tmp[1687]*kernel[8];
				ans[1587]<=tmp[1486]*kernel[0]+tmp[1487]*kernel[1]+tmp[1488]*kernel[2]+tmp[1586]*kernel[3]+tmp[1587]*kernel[4]+tmp[1588]*kernel[5]+tmp[1686]*kernel[6]+tmp[1687]*kernel[7]+tmp[1688]*kernel[8];
				ans[1588]<=tmp[1487]*kernel[0]+tmp[1488]*kernel[1]+tmp[1489]*kernel[2]+tmp[1587]*kernel[3]+tmp[1588]*kernel[4]+tmp[1589]*kernel[5]+tmp[1687]*kernel[6]+tmp[1688]*kernel[7]+tmp[1689]*kernel[8];
				ans[1589]<=tmp[1488]*kernel[0]+tmp[1489]*kernel[1]+tmp[1490]*kernel[2]+tmp[1588]*kernel[3]+tmp[1589]*kernel[4]+tmp[1590]*kernel[5]+tmp[1688]*kernel[6]+tmp[1689]*kernel[7]+tmp[1690]*kernel[8];
				ans[1590]<=tmp[1489]*kernel[0]+tmp[1490]*kernel[1]+tmp[1491]*kernel[2]+tmp[1589]*kernel[3]+tmp[1590]*kernel[4]+tmp[1591]*kernel[5]+tmp[1689]*kernel[6]+tmp[1690]*kernel[7]+tmp[1691]*kernel[8];
				ans[1591]<=tmp[1490]*kernel[0]+tmp[1491]*kernel[1]+tmp[1492]*kernel[2]+tmp[1590]*kernel[3]+tmp[1591]*kernel[4]+tmp[1592]*kernel[5]+tmp[1690]*kernel[6]+tmp[1691]*kernel[7]+tmp[1692]*kernel[8];
				ans[1592]<=tmp[1491]*kernel[0]+tmp[1492]*kernel[1]+tmp[1493]*kernel[2]+tmp[1591]*kernel[3]+tmp[1592]*kernel[4]+tmp[1593]*kernel[5]+tmp[1691]*kernel[6]+tmp[1692]*kernel[7]+tmp[1693]*kernel[8];
				ans[1593]<=tmp[1492]*kernel[0]+tmp[1493]*kernel[1]+tmp[1494]*kernel[2]+tmp[1592]*kernel[3]+tmp[1593]*kernel[4]+tmp[1594]*kernel[5]+tmp[1692]*kernel[6]+tmp[1693]*kernel[7]+tmp[1694]*kernel[8];
				ans[1594]<=tmp[1493]*kernel[0]+tmp[1494]*kernel[1]+tmp[1495]*kernel[2]+tmp[1593]*kernel[3]+tmp[1594]*kernel[4]+tmp[1595]*kernel[5]+tmp[1693]*kernel[6]+tmp[1694]*kernel[7]+tmp[1695]*kernel[8];
				ans[1595]<=tmp[1494]*kernel[0]+tmp[1495]*kernel[1]+tmp[1496]*kernel[2]+tmp[1594]*kernel[3]+tmp[1595]*kernel[4]+tmp[1596]*kernel[5]+tmp[1694]*kernel[6]+tmp[1695]*kernel[7]+tmp[1696]*kernel[8];
				ans[1596]<=tmp[1495]*kernel[0]+tmp[1496]*kernel[1]+tmp[1497]*kernel[2]+tmp[1595]*kernel[3]+tmp[1596]*kernel[4]+tmp[1597]*kernel[5]+tmp[1695]*kernel[6]+tmp[1696]*kernel[7]+tmp[1697]*kernel[8];
				ans[1597]<=tmp[1496]*kernel[0]+tmp[1497]*kernel[1]+tmp[1498]*kernel[2]+tmp[1596]*kernel[3]+tmp[1597]*kernel[4]+tmp[1598]*kernel[5]+tmp[1696]*kernel[6]+tmp[1697]*kernel[7]+tmp[1698]*kernel[8];
				ans[1598]<=tmp[1497]*kernel[0]+tmp[1498]*kernel[1]+tmp[1499]*kernel[2]+tmp[1597]*kernel[3]+tmp[1598]*kernel[4]+tmp[1599]*kernel[5]+tmp[1697]*kernel[6]+tmp[1698]*kernel[7]+tmp[1699]*kernel[8];
				ans[1599]<=tmp[1498]*kernel[0]+tmp[1499]*kernel[1]+tmp[1598]*kernel[3]+tmp[1599]*kernel[4]+tmp[1698]*kernel[6]+tmp[1699]*kernel[7];
				ans[1600]<=tmp[1500]*kernel[1]+tmp[1501]*kernel[2]+tmp[1600]*kernel[4]+tmp[1601]*kernel[5]+tmp[1700]*kernel[7]+tmp[1701]*kernel[8];
				ans[1601]<=tmp[1500]*kernel[0]+tmp[1501]*kernel[1]+tmp[1502]*kernel[2]+tmp[1600]*kernel[3]+tmp[1601]*kernel[4]+tmp[1602]*kernel[5]+tmp[1700]*kernel[6]+tmp[1701]*kernel[7]+tmp[1702]*kernel[8];
				ans[1602]<=tmp[1501]*kernel[0]+tmp[1502]*kernel[1]+tmp[1503]*kernel[2]+tmp[1601]*kernel[3]+tmp[1602]*kernel[4]+tmp[1603]*kernel[5]+tmp[1701]*kernel[6]+tmp[1702]*kernel[7]+tmp[1703]*kernel[8];
				ans[1603]<=tmp[1502]*kernel[0]+tmp[1503]*kernel[1]+tmp[1504]*kernel[2]+tmp[1602]*kernel[3]+tmp[1603]*kernel[4]+tmp[1604]*kernel[5]+tmp[1702]*kernel[6]+tmp[1703]*kernel[7]+tmp[1704]*kernel[8];
				ans[1604]<=tmp[1503]*kernel[0]+tmp[1504]*kernel[1]+tmp[1505]*kernel[2]+tmp[1603]*kernel[3]+tmp[1604]*kernel[4]+tmp[1605]*kernel[5]+tmp[1703]*kernel[6]+tmp[1704]*kernel[7]+tmp[1705]*kernel[8];
				ans[1605]<=tmp[1504]*kernel[0]+tmp[1505]*kernel[1]+tmp[1506]*kernel[2]+tmp[1604]*kernel[3]+tmp[1605]*kernel[4]+tmp[1606]*kernel[5]+tmp[1704]*kernel[6]+tmp[1705]*kernel[7]+tmp[1706]*kernel[8];
				ans[1606]<=tmp[1505]*kernel[0]+tmp[1506]*kernel[1]+tmp[1507]*kernel[2]+tmp[1605]*kernel[3]+tmp[1606]*kernel[4]+tmp[1607]*kernel[5]+tmp[1705]*kernel[6]+tmp[1706]*kernel[7]+tmp[1707]*kernel[8];
				ans[1607]<=tmp[1506]*kernel[0]+tmp[1507]*kernel[1]+tmp[1508]*kernel[2]+tmp[1606]*kernel[3]+tmp[1607]*kernel[4]+tmp[1608]*kernel[5]+tmp[1706]*kernel[6]+tmp[1707]*kernel[7]+tmp[1708]*kernel[8];
				ans[1608]<=tmp[1507]*kernel[0]+tmp[1508]*kernel[1]+tmp[1509]*kernel[2]+tmp[1607]*kernel[3]+tmp[1608]*kernel[4]+tmp[1609]*kernel[5]+tmp[1707]*kernel[6]+tmp[1708]*kernel[7]+tmp[1709]*kernel[8];
				ans[1609]<=tmp[1508]*kernel[0]+tmp[1509]*kernel[1]+tmp[1510]*kernel[2]+tmp[1608]*kernel[3]+tmp[1609]*kernel[4]+tmp[1610]*kernel[5]+tmp[1708]*kernel[6]+tmp[1709]*kernel[7]+tmp[1710]*kernel[8];
				ans[1610]<=tmp[1509]*kernel[0]+tmp[1510]*kernel[1]+tmp[1511]*kernel[2]+tmp[1609]*kernel[3]+tmp[1610]*kernel[4]+tmp[1611]*kernel[5]+tmp[1709]*kernel[6]+tmp[1710]*kernel[7]+tmp[1711]*kernel[8];
				ans[1611]<=tmp[1510]*kernel[0]+tmp[1511]*kernel[1]+tmp[1512]*kernel[2]+tmp[1610]*kernel[3]+tmp[1611]*kernel[4]+tmp[1612]*kernel[5]+tmp[1710]*kernel[6]+tmp[1711]*kernel[7]+tmp[1712]*kernel[8];
				ans[1612]<=tmp[1511]*kernel[0]+tmp[1512]*kernel[1]+tmp[1513]*kernel[2]+tmp[1611]*kernel[3]+tmp[1612]*kernel[4]+tmp[1613]*kernel[5]+tmp[1711]*kernel[6]+tmp[1712]*kernel[7]+tmp[1713]*kernel[8];
				ans[1613]<=tmp[1512]*kernel[0]+tmp[1513]*kernel[1]+tmp[1514]*kernel[2]+tmp[1612]*kernel[3]+tmp[1613]*kernel[4]+tmp[1614]*kernel[5]+tmp[1712]*kernel[6]+tmp[1713]*kernel[7]+tmp[1714]*kernel[8];
				ans[1614]<=tmp[1513]*kernel[0]+tmp[1514]*kernel[1]+tmp[1515]*kernel[2]+tmp[1613]*kernel[3]+tmp[1614]*kernel[4]+tmp[1615]*kernel[5]+tmp[1713]*kernel[6]+tmp[1714]*kernel[7]+tmp[1715]*kernel[8];
				ans[1615]<=tmp[1514]*kernel[0]+tmp[1515]*kernel[1]+tmp[1516]*kernel[2]+tmp[1614]*kernel[3]+tmp[1615]*kernel[4]+tmp[1616]*kernel[5]+tmp[1714]*kernel[6]+tmp[1715]*kernel[7]+tmp[1716]*kernel[8];
				ans[1616]<=tmp[1515]*kernel[0]+tmp[1516]*kernel[1]+tmp[1517]*kernel[2]+tmp[1615]*kernel[3]+tmp[1616]*kernel[4]+tmp[1617]*kernel[5]+tmp[1715]*kernel[6]+tmp[1716]*kernel[7]+tmp[1717]*kernel[8];
				ans[1617]<=tmp[1516]*kernel[0]+tmp[1517]*kernel[1]+tmp[1518]*kernel[2]+tmp[1616]*kernel[3]+tmp[1617]*kernel[4]+tmp[1618]*kernel[5]+tmp[1716]*kernel[6]+tmp[1717]*kernel[7]+tmp[1718]*kernel[8];
				ans[1618]<=tmp[1517]*kernel[0]+tmp[1518]*kernel[1]+tmp[1519]*kernel[2]+tmp[1617]*kernel[3]+tmp[1618]*kernel[4]+tmp[1619]*kernel[5]+tmp[1717]*kernel[6]+tmp[1718]*kernel[7]+tmp[1719]*kernel[8];
				ans[1619]<=tmp[1518]*kernel[0]+tmp[1519]*kernel[1]+tmp[1520]*kernel[2]+tmp[1618]*kernel[3]+tmp[1619]*kernel[4]+tmp[1620]*kernel[5]+tmp[1718]*kernel[6]+tmp[1719]*kernel[7]+tmp[1720]*kernel[8];
				ans[1620]<=tmp[1519]*kernel[0]+tmp[1520]*kernel[1]+tmp[1521]*kernel[2]+tmp[1619]*kernel[3]+tmp[1620]*kernel[4]+tmp[1621]*kernel[5]+tmp[1719]*kernel[6]+tmp[1720]*kernel[7]+tmp[1721]*kernel[8];
				ans[1621]<=tmp[1520]*kernel[0]+tmp[1521]*kernel[1]+tmp[1522]*kernel[2]+tmp[1620]*kernel[3]+tmp[1621]*kernel[4]+tmp[1622]*kernel[5]+tmp[1720]*kernel[6]+tmp[1721]*kernel[7]+tmp[1722]*kernel[8];
				ans[1622]<=tmp[1521]*kernel[0]+tmp[1522]*kernel[1]+tmp[1523]*kernel[2]+tmp[1621]*kernel[3]+tmp[1622]*kernel[4]+tmp[1623]*kernel[5]+tmp[1721]*kernel[6]+tmp[1722]*kernel[7]+tmp[1723]*kernel[8];
				ans[1623]<=tmp[1522]*kernel[0]+tmp[1523]*kernel[1]+tmp[1524]*kernel[2]+tmp[1622]*kernel[3]+tmp[1623]*kernel[4]+tmp[1624]*kernel[5]+tmp[1722]*kernel[6]+tmp[1723]*kernel[7]+tmp[1724]*kernel[8];
				ans[1624]<=tmp[1523]*kernel[0]+tmp[1524]*kernel[1]+tmp[1525]*kernel[2]+tmp[1623]*kernel[3]+tmp[1624]*kernel[4]+tmp[1625]*kernel[5]+tmp[1723]*kernel[6]+tmp[1724]*kernel[7]+tmp[1725]*kernel[8];
				ans[1625]<=tmp[1524]*kernel[0]+tmp[1525]*kernel[1]+tmp[1526]*kernel[2]+tmp[1624]*kernel[3]+tmp[1625]*kernel[4]+tmp[1626]*kernel[5]+tmp[1724]*kernel[6]+tmp[1725]*kernel[7]+tmp[1726]*kernel[8];
				ans[1626]<=tmp[1525]*kernel[0]+tmp[1526]*kernel[1]+tmp[1527]*kernel[2]+tmp[1625]*kernel[3]+tmp[1626]*kernel[4]+tmp[1627]*kernel[5]+tmp[1725]*kernel[6]+tmp[1726]*kernel[7]+tmp[1727]*kernel[8];
				ans[1627]<=tmp[1526]*kernel[0]+tmp[1527]*kernel[1]+tmp[1528]*kernel[2]+tmp[1626]*kernel[3]+tmp[1627]*kernel[4]+tmp[1628]*kernel[5]+tmp[1726]*kernel[6]+tmp[1727]*kernel[7]+tmp[1728]*kernel[8];
				ans[1628]<=tmp[1527]*kernel[0]+tmp[1528]*kernel[1]+tmp[1529]*kernel[2]+tmp[1627]*kernel[3]+tmp[1628]*kernel[4]+tmp[1629]*kernel[5]+tmp[1727]*kernel[6]+tmp[1728]*kernel[7]+tmp[1729]*kernel[8];
				ans[1629]<=tmp[1528]*kernel[0]+tmp[1529]*kernel[1]+tmp[1530]*kernel[2]+tmp[1628]*kernel[3]+tmp[1629]*kernel[4]+tmp[1630]*kernel[5]+tmp[1728]*kernel[6]+tmp[1729]*kernel[7]+tmp[1730]*kernel[8];
				ans[1630]<=tmp[1529]*kernel[0]+tmp[1530]*kernel[1]+tmp[1531]*kernel[2]+tmp[1629]*kernel[3]+tmp[1630]*kernel[4]+tmp[1631]*kernel[5]+tmp[1729]*kernel[6]+tmp[1730]*kernel[7]+tmp[1731]*kernel[8];
				ans[1631]<=tmp[1530]*kernel[0]+tmp[1531]*kernel[1]+tmp[1532]*kernel[2]+tmp[1630]*kernel[3]+tmp[1631]*kernel[4]+tmp[1632]*kernel[5]+tmp[1730]*kernel[6]+tmp[1731]*kernel[7]+tmp[1732]*kernel[8];
				ans[1632]<=tmp[1531]*kernel[0]+tmp[1532]*kernel[1]+tmp[1533]*kernel[2]+tmp[1631]*kernel[3]+tmp[1632]*kernel[4]+tmp[1633]*kernel[5]+tmp[1731]*kernel[6]+tmp[1732]*kernel[7]+tmp[1733]*kernel[8];
				ans[1633]<=tmp[1532]*kernel[0]+tmp[1533]*kernel[1]+tmp[1534]*kernel[2]+tmp[1632]*kernel[3]+tmp[1633]*kernel[4]+tmp[1634]*kernel[5]+tmp[1732]*kernel[6]+tmp[1733]*kernel[7]+tmp[1734]*kernel[8];
				ans[1634]<=tmp[1533]*kernel[0]+tmp[1534]*kernel[1]+tmp[1535]*kernel[2]+tmp[1633]*kernel[3]+tmp[1634]*kernel[4]+tmp[1635]*kernel[5]+tmp[1733]*kernel[6]+tmp[1734]*kernel[7]+tmp[1735]*kernel[8];
				ans[1635]<=tmp[1534]*kernel[0]+tmp[1535]*kernel[1]+tmp[1536]*kernel[2]+tmp[1634]*kernel[3]+tmp[1635]*kernel[4]+tmp[1636]*kernel[5]+tmp[1734]*kernel[6]+tmp[1735]*kernel[7]+tmp[1736]*kernel[8];
				ans[1636]<=tmp[1535]*kernel[0]+tmp[1536]*kernel[1]+tmp[1537]*kernel[2]+tmp[1635]*kernel[3]+tmp[1636]*kernel[4]+tmp[1637]*kernel[5]+tmp[1735]*kernel[6]+tmp[1736]*kernel[7]+tmp[1737]*kernel[8];
				ans[1637]<=tmp[1536]*kernel[0]+tmp[1537]*kernel[1]+tmp[1538]*kernel[2]+tmp[1636]*kernel[3]+tmp[1637]*kernel[4]+tmp[1638]*kernel[5]+tmp[1736]*kernel[6]+tmp[1737]*kernel[7]+tmp[1738]*kernel[8];
				ans[1638]<=tmp[1537]*kernel[0]+tmp[1538]*kernel[1]+tmp[1539]*kernel[2]+tmp[1637]*kernel[3]+tmp[1638]*kernel[4]+tmp[1639]*kernel[5]+tmp[1737]*kernel[6]+tmp[1738]*kernel[7]+tmp[1739]*kernel[8];
				ans[1639]<=tmp[1538]*kernel[0]+tmp[1539]*kernel[1]+tmp[1540]*kernel[2]+tmp[1638]*kernel[3]+tmp[1639]*kernel[4]+tmp[1640]*kernel[5]+tmp[1738]*kernel[6]+tmp[1739]*kernel[7]+tmp[1740]*kernel[8];
				ans[1640]<=tmp[1539]*kernel[0]+tmp[1540]*kernel[1]+tmp[1541]*kernel[2]+tmp[1639]*kernel[3]+tmp[1640]*kernel[4]+tmp[1641]*kernel[5]+tmp[1739]*kernel[6]+tmp[1740]*kernel[7]+tmp[1741]*kernel[8];
				ans[1641]<=tmp[1540]*kernel[0]+tmp[1541]*kernel[1]+tmp[1542]*kernel[2]+tmp[1640]*kernel[3]+tmp[1641]*kernel[4]+tmp[1642]*kernel[5]+tmp[1740]*kernel[6]+tmp[1741]*kernel[7]+tmp[1742]*kernel[8];
				ans[1642]<=tmp[1541]*kernel[0]+tmp[1542]*kernel[1]+tmp[1543]*kernel[2]+tmp[1641]*kernel[3]+tmp[1642]*kernel[4]+tmp[1643]*kernel[5]+tmp[1741]*kernel[6]+tmp[1742]*kernel[7]+tmp[1743]*kernel[8];
				ans[1643]<=tmp[1542]*kernel[0]+tmp[1543]*kernel[1]+tmp[1544]*kernel[2]+tmp[1642]*kernel[3]+tmp[1643]*kernel[4]+tmp[1644]*kernel[5]+tmp[1742]*kernel[6]+tmp[1743]*kernel[7]+tmp[1744]*kernel[8];
				ans[1644]<=tmp[1543]*kernel[0]+tmp[1544]*kernel[1]+tmp[1545]*kernel[2]+tmp[1643]*kernel[3]+tmp[1644]*kernel[4]+tmp[1645]*kernel[5]+tmp[1743]*kernel[6]+tmp[1744]*kernel[7]+tmp[1745]*kernel[8];
				ans[1645]<=tmp[1544]*kernel[0]+tmp[1545]*kernel[1]+tmp[1546]*kernel[2]+tmp[1644]*kernel[3]+tmp[1645]*kernel[4]+tmp[1646]*kernel[5]+tmp[1744]*kernel[6]+tmp[1745]*kernel[7]+tmp[1746]*kernel[8];
				ans[1646]<=tmp[1545]*kernel[0]+tmp[1546]*kernel[1]+tmp[1547]*kernel[2]+tmp[1645]*kernel[3]+tmp[1646]*kernel[4]+tmp[1647]*kernel[5]+tmp[1745]*kernel[6]+tmp[1746]*kernel[7]+tmp[1747]*kernel[8];
				ans[1647]<=tmp[1546]*kernel[0]+tmp[1547]*kernel[1]+tmp[1548]*kernel[2]+tmp[1646]*kernel[3]+tmp[1647]*kernel[4]+tmp[1648]*kernel[5]+tmp[1746]*kernel[6]+tmp[1747]*kernel[7]+tmp[1748]*kernel[8];
				ans[1648]<=tmp[1547]*kernel[0]+tmp[1548]*kernel[1]+tmp[1549]*kernel[2]+tmp[1647]*kernel[3]+tmp[1648]*kernel[4]+tmp[1649]*kernel[5]+tmp[1747]*kernel[6]+tmp[1748]*kernel[7]+tmp[1749]*kernel[8];
				ans[1649]<=tmp[1548]*kernel[0]+tmp[1549]*kernel[1]+tmp[1550]*kernel[2]+tmp[1648]*kernel[3]+tmp[1649]*kernel[4]+tmp[1650]*kernel[5]+tmp[1748]*kernel[6]+tmp[1749]*kernel[7]+tmp[1750]*kernel[8];
				ans[1650]<=tmp[1549]*kernel[0]+tmp[1550]*kernel[1]+tmp[1551]*kernel[2]+tmp[1649]*kernel[3]+tmp[1650]*kernel[4]+tmp[1651]*kernel[5]+tmp[1749]*kernel[6]+tmp[1750]*kernel[7]+tmp[1751]*kernel[8];
				ans[1651]<=tmp[1550]*kernel[0]+tmp[1551]*kernel[1]+tmp[1552]*kernel[2]+tmp[1650]*kernel[3]+tmp[1651]*kernel[4]+tmp[1652]*kernel[5]+tmp[1750]*kernel[6]+tmp[1751]*kernel[7]+tmp[1752]*kernel[8];
				ans[1652]<=tmp[1551]*kernel[0]+tmp[1552]*kernel[1]+tmp[1553]*kernel[2]+tmp[1651]*kernel[3]+tmp[1652]*kernel[4]+tmp[1653]*kernel[5]+tmp[1751]*kernel[6]+tmp[1752]*kernel[7]+tmp[1753]*kernel[8];
				ans[1653]<=tmp[1552]*kernel[0]+tmp[1553]*kernel[1]+tmp[1554]*kernel[2]+tmp[1652]*kernel[3]+tmp[1653]*kernel[4]+tmp[1654]*kernel[5]+tmp[1752]*kernel[6]+tmp[1753]*kernel[7]+tmp[1754]*kernel[8];
				ans[1654]<=tmp[1553]*kernel[0]+tmp[1554]*kernel[1]+tmp[1555]*kernel[2]+tmp[1653]*kernel[3]+tmp[1654]*kernel[4]+tmp[1655]*kernel[5]+tmp[1753]*kernel[6]+tmp[1754]*kernel[7]+tmp[1755]*kernel[8];
				ans[1655]<=tmp[1554]*kernel[0]+tmp[1555]*kernel[1]+tmp[1556]*kernel[2]+tmp[1654]*kernel[3]+tmp[1655]*kernel[4]+tmp[1656]*kernel[5]+tmp[1754]*kernel[6]+tmp[1755]*kernel[7]+tmp[1756]*kernel[8];
				ans[1656]<=tmp[1555]*kernel[0]+tmp[1556]*kernel[1]+tmp[1557]*kernel[2]+tmp[1655]*kernel[3]+tmp[1656]*kernel[4]+tmp[1657]*kernel[5]+tmp[1755]*kernel[6]+tmp[1756]*kernel[7]+tmp[1757]*kernel[8];
				ans[1657]<=tmp[1556]*kernel[0]+tmp[1557]*kernel[1]+tmp[1558]*kernel[2]+tmp[1656]*kernel[3]+tmp[1657]*kernel[4]+tmp[1658]*kernel[5]+tmp[1756]*kernel[6]+tmp[1757]*kernel[7]+tmp[1758]*kernel[8];
				ans[1658]<=tmp[1557]*kernel[0]+tmp[1558]*kernel[1]+tmp[1559]*kernel[2]+tmp[1657]*kernel[3]+tmp[1658]*kernel[4]+tmp[1659]*kernel[5]+tmp[1757]*kernel[6]+tmp[1758]*kernel[7]+tmp[1759]*kernel[8];
				ans[1659]<=tmp[1558]*kernel[0]+tmp[1559]*kernel[1]+tmp[1560]*kernel[2]+tmp[1658]*kernel[3]+tmp[1659]*kernel[4]+tmp[1660]*kernel[5]+tmp[1758]*kernel[6]+tmp[1759]*kernel[7]+tmp[1760]*kernel[8];
				ans[1660]<=tmp[1559]*kernel[0]+tmp[1560]*kernel[1]+tmp[1561]*kernel[2]+tmp[1659]*kernel[3]+tmp[1660]*kernel[4]+tmp[1661]*kernel[5]+tmp[1759]*kernel[6]+tmp[1760]*kernel[7]+tmp[1761]*kernel[8];
				ans[1661]<=tmp[1560]*kernel[0]+tmp[1561]*kernel[1]+tmp[1562]*kernel[2]+tmp[1660]*kernel[3]+tmp[1661]*kernel[4]+tmp[1662]*kernel[5]+tmp[1760]*kernel[6]+tmp[1761]*kernel[7]+tmp[1762]*kernel[8];
				ans[1662]<=tmp[1561]*kernel[0]+tmp[1562]*kernel[1]+tmp[1563]*kernel[2]+tmp[1661]*kernel[3]+tmp[1662]*kernel[4]+tmp[1663]*kernel[5]+tmp[1761]*kernel[6]+tmp[1762]*kernel[7]+tmp[1763]*kernel[8];
				ans[1663]<=tmp[1562]*kernel[0]+tmp[1563]*kernel[1]+tmp[1564]*kernel[2]+tmp[1662]*kernel[3]+tmp[1663]*kernel[4]+tmp[1664]*kernel[5]+tmp[1762]*kernel[6]+tmp[1763]*kernel[7]+tmp[1764]*kernel[8];
				ans[1664]<=tmp[1563]*kernel[0]+tmp[1564]*kernel[1]+tmp[1565]*kernel[2]+tmp[1663]*kernel[3]+tmp[1664]*kernel[4]+tmp[1665]*kernel[5]+tmp[1763]*kernel[6]+tmp[1764]*kernel[7]+tmp[1765]*kernel[8];
				ans[1665]<=tmp[1564]*kernel[0]+tmp[1565]*kernel[1]+tmp[1566]*kernel[2]+tmp[1664]*kernel[3]+tmp[1665]*kernel[4]+tmp[1666]*kernel[5]+tmp[1764]*kernel[6]+tmp[1765]*kernel[7]+tmp[1766]*kernel[8];
				ans[1666]<=tmp[1565]*kernel[0]+tmp[1566]*kernel[1]+tmp[1567]*kernel[2]+tmp[1665]*kernel[3]+tmp[1666]*kernel[4]+tmp[1667]*kernel[5]+tmp[1765]*kernel[6]+tmp[1766]*kernel[7]+tmp[1767]*kernel[8];
				ans[1667]<=tmp[1566]*kernel[0]+tmp[1567]*kernel[1]+tmp[1568]*kernel[2]+tmp[1666]*kernel[3]+tmp[1667]*kernel[4]+tmp[1668]*kernel[5]+tmp[1766]*kernel[6]+tmp[1767]*kernel[7]+tmp[1768]*kernel[8];
				ans[1668]<=tmp[1567]*kernel[0]+tmp[1568]*kernel[1]+tmp[1569]*kernel[2]+tmp[1667]*kernel[3]+tmp[1668]*kernel[4]+tmp[1669]*kernel[5]+tmp[1767]*kernel[6]+tmp[1768]*kernel[7]+tmp[1769]*kernel[8];
				ans[1669]<=tmp[1568]*kernel[0]+tmp[1569]*kernel[1]+tmp[1570]*kernel[2]+tmp[1668]*kernel[3]+tmp[1669]*kernel[4]+tmp[1670]*kernel[5]+tmp[1768]*kernel[6]+tmp[1769]*kernel[7]+tmp[1770]*kernel[8];
				ans[1670]<=tmp[1569]*kernel[0]+tmp[1570]*kernel[1]+tmp[1571]*kernel[2]+tmp[1669]*kernel[3]+tmp[1670]*kernel[4]+tmp[1671]*kernel[5]+tmp[1769]*kernel[6]+tmp[1770]*kernel[7]+tmp[1771]*kernel[8];
				ans[1671]<=tmp[1570]*kernel[0]+tmp[1571]*kernel[1]+tmp[1572]*kernel[2]+tmp[1670]*kernel[3]+tmp[1671]*kernel[4]+tmp[1672]*kernel[5]+tmp[1770]*kernel[6]+tmp[1771]*kernel[7]+tmp[1772]*kernel[8];
				ans[1672]<=tmp[1571]*kernel[0]+tmp[1572]*kernel[1]+tmp[1573]*kernel[2]+tmp[1671]*kernel[3]+tmp[1672]*kernel[4]+tmp[1673]*kernel[5]+tmp[1771]*kernel[6]+tmp[1772]*kernel[7]+tmp[1773]*kernel[8];
				ans[1673]<=tmp[1572]*kernel[0]+tmp[1573]*kernel[1]+tmp[1574]*kernel[2]+tmp[1672]*kernel[3]+tmp[1673]*kernel[4]+tmp[1674]*kernel[5]+tmp[1772]*kernel[6]+tmp[1773]*kernel[7]+tmp[1774]*kernel[8];
				ans[1674]<=tmp[1573]*kernel[0]+tmp[1574]*kernel[1]+tmp[1575]*kernel[2]+tmp[1673]*kernel[3]+tmp[1674]*kernel[4]+tmp[1675]*kernel[5]+tmp[1773]*kernel[6]+tmp[1774]*kernel[7]+tmp[1775]*kernel[8];
				ans[1675]<=tmp[1574]*kernel[0]+tmp[1575]*kernel[1]+tmp[1576]*kernel[2]+tmp[1674]*kernel[3]+tmp[1675]*kernel[4]+tmp[1676]*kernel[5]+tmp[1774]*kernel[6]+tmp[1775]*kernel[7]+tmp[1776]*kernel[8];
				ans[1676]<=tmp[1575]*kernel[0]+tmp[1576]*kernel[1]+tmp[1577]*kernel[2]+tmp[1675]*kernel[3]+tmp[1676]*kernel[4]+tmp[1677]*kernel[5]+tmp[1775]*kernel[6]+tmp[1776]*kernel[7]+tmp[1777]*kernel[8];
				ans[1677]<=tmp[1576]*kernel[0]+tmp[1577]*kernel[1]+tmp[1578]*kernel[2]+tmp[1676]*kernel[3]+tmp[1677]*kernel[4]+tmp[1678]*kernel[5]+tmp[1776]*kernel[6]+tmp[1777]*kernel[7]+tmp[1778]*kernel[8];
				ans[1678]<=tmp[1577]*kernel[0]+tmp[1578]*kernel[1]+tmp[1579]*kernel[2]+tmp[1677]*kernel[3]+tmp[1678]*kernel[4]+tmp[1679]*kernel[5]+tmp[1777]*kernel[6]+tmp[1778]*kernel[7]+tmp[1779]*kernel[8];
				ans[1679]<=tmp[1578]*kernel[0]+tmp[1579]*kernel[1]+tmp[1580]*kernel[2]+tmp[1678]*kernel[3]+tmp[1679]*kernel[4]+tmp[1680]*kernel[5]+tmp[1778]*kernel[6]+tmp[1779]*kernel[7]+tmp[1780]*kernel[8];
				ans[1680]<=tmp[1579]*kernel[0]+tmp[1580]*kernel[1]+tmp[1581]*kernel[2]+tmp[1679]*kernel[3]+tmp[1680]*kernel[4]+tmp[1681]*kernel[5]+tmp[1779]*kernel[6]+tmp[1780]*kernel[7]+tmp[1781]*kernel[8];
				ans[1681]<=tmp[1580]*kernel[0]+tmp[1581]*kernel[1]+tmp[1582]*kernel[2]+tmp[1680]*kernel[3]+tmp[1681]*kernel[4]+tmp[1682]*kernel[5]+tmp[1780]*kernel[6]+tmp[1781]*kernel[7]+tmp[1782]*kernel[8];
				ans[1682]<=tmp[1581]*kernel[0]+tmp[1582]*kernel[1]+tmp[1583]*kernel[2]+tmp[1681]*kernel[3]+tmp[1682]*kernel[4]+tmp[1683]*kernel[5]+tmp[1781]*kernel[6]+tmp[1782]*kernel[7]+tmp[1783]*kernel[8];
				ans[1683]<=tmp[1582]*kernel[0]+tmp[1583]*kernel[1]+tmp[1584]*kernel[2]+tmp[1682]*kernel[3]+tmp[1683]*kernel[4]+tmp[1684]*kernel[5]+tmp[1782]*kernel[6]+tmp[1783]*kernel[7]+tmp[1784]*kernel[8];
				ans[1684]<=tmp[1583]*kernel[0]+tmp[1584]*kernel[1]+tmp[1585]*kernel[2]+tmp[1683]*kernel[3]+tmp[1684]*kernel[4]+tmp[1685]*kernel[5]+tmp[1783]*kernel[6]+tmp[1784]*kernel[7]+tmp[1785]*kernel[8];
				ans[1685]<=tmp[1584]*kernel[0]+tmp[1585]*kernel[1]+tmp[1586]*kernel[2]+tmp[1684]*kernel[3]+tmp[1685]*kernel[4]+tmp[1686]*kernel[5]+tmp[1784]*kernel[6]+tmp[1785]*kernel[7]+tmp[1786]*kernel[8];
				ans[1686]<=tmp[1585]*kernel[0]+tmp[1586]*kernel[1]+tmp[1587]*kernel[2]+tmp[1685]*kernel[3]+tmp[1686]*kernel[4]+tmp[1687]*kernel[5]+tmp[1785]*kernel[6]+tmp[1786]*kernel[7]+tmp[1787]*kernel[8];
				ans[1687]<=tmp[1586]*kernel[0]+tmp[1587]*kernel[1]+tmp[1588]*kernel[2]+tmp[1686]*kernel[3]+tmp[1687]*kernel[4]+tmp[1688]*kernel[5]+tmp[1786]*kernel[6]+tmp[1787]*kernel[7]+tmp[1788]*kernel[8];
				ans[1688]<=tmp[1587]*kernel[0]+tmp[1588]*kernel[1]+tmp[1589]*kernel[2]+tmp[1687]*kernel[3]+tmp[1688]*kernel[4]+tmp[1689]*kernel[5]+tmp[1787]*kernel[6]+tmp[1788]*kernel[7]+tmp[1789]*kernel[8];
				ans[1689]<=tmp[1588]*kernel[0]+tmp[1589]*kernel[1]+tmp[1590]*kernel[2]+tmp[1688]*kernel[3]+tmp[1689]*kernel[4]+tmp[1690]*kernel[5]+tmp[1788]*kernel[6]+tmp[1789]*kernel[7]+tmp[1790]*kernel[8];
				ans[1690]<=tmp[1589]*kernel[0]+tmp[1590]*kernel[1]+tmp[1591]*kernel[2]+tmp[1689]*kernel[3]+tmp[1690]*kernel[4]+tmp[1691]*kernel[5]+tmp[1789]*kernel[6]+tmp[1790]*kernel[7]+tmp[1791]*kernel[8];
				ans[1691]<=tmp[1590]*kernel[0]+tmp[1591]*kernel[1]+tmp[1592]*kernel[2]+tmp[1690]*kernel[3]+tmp[1691]*kernel[4]+tmp[1692]*kernel[5]+tmp[1790]*kernel[6]+tmp[1791]*kernel[7]+tmp[1792]*kernel[8];
				ans[1692]<=tmp[1591]*kernel[0]+tmp[1592]*kernel[1]+tmp[1593]*kernel[2]+tmp[1691]*kernel[3]+tmp[1692]*kernel[4]+tmp[1693]*kernel[5]+tmp[1791]*kernel[6]+tmp[1792]*kernel[7]+tmp[1793]*kernel[8];
				ans[1693]<=tmp[1592]*kernel[0]+tmp[1593]*kernel[1]+tmp[1594]*kernel[2]+tmp[1692]*kernel[3]+tmp[1693]*kernel[4]+tmp[1694]*kernel[5]+tmp[1792]*kernel[6]+tmp[1793]*kernel[7]+tmp[1794]*kernel[8];
				ans[1694]<=tmp[1593]*kernel[0]+tmp[1594]*kernel[1]+tmp[1595]*kernel[2]+tmp[1693]*kernel[3]+tmp[1694]*kernel[4]+tmp[1695]*kernel[5]+tmp[1793]*kernel[6]+tmp[1794]*kernel[7]+tmp[1795]*kernel[8];
				ans[1695]<=tmp[1594]*kernel[0]+tmp[1595]*kernel[1]+tmp[1596]*kernel[2]+tmp[1694]*kernel[3]+tmp[1695]*kernel[4]+tmp[1696]*kernel[5]+tmp[1794]*kernel[6]+tmp[1795]*kernel[7]+tmp[1796]*kernel[8];
				ans[1696]<=tmp[1595]*kernel[0]+tmp[1596]*kernel[1]+tmp[1597]*kernel[2]+tmp[1695]*kernel[3]+tmp[1696]*kernel[4]+tmp[1697]*kernel[5]+tmp[1795]*kernel[6]+tmp[1796]*kernel[7]+tmp[1797]*kernel[8];
				ans[1697]<=tmp[1596]*kernel[0]+tmp[1597]*kernel[1]+tmp[1598]*kernel[2]+tmp[1696]*kernel[3]+tmp[1697]*kernel[4]+tmp[1698]*kernel[5]+tmp[1796]*kernel[6]+tmp[1797]*kernel[7]+tmp[1798]*kernel[8];
				ans[1698]<=tmp[1597]*kernel[0]+tmp[1598]*kernel[1]+tmp[1599]*kernel[2]+tmp[1697]*kernel[3]+tmp[1698]*kernel[4]+tmp[1699]*kernel[5]+tmp[1797]*kernel[6]+tmp[1798]*kernel[7]+tmp[1799]*kernel[8];
				ans[1699]<=tmp[1598]*kernel[0]+tmp[1599]*kernel[1]+tmp[1698]*kernel[3]+tmp[1699]*kernel[4]+tmp[1798]*kernel[6]+tmp[1799]*kernel[7];
				ans[1700]<=tmp[1600]*kernel[1]+tmp[1601]*kernel[2]+tmp[1700]*kernel[4]+tmp[1701]*kernel[5]+tmp[1800]*kernel[7]+tmp[1801]*kernel[8];
				ans[1701]<=tmp[1600]*kernel[0]+tmp[1601]*kernel[1]+tmp[1602]*kernel[2]+tmp[1700]*kernel[3]+tmp[1701]*kernel[4]+tmp[1702]*kernel[5]+tmp[1800]*kernel[6]+tmp[1801]*kernel[7]+tmp[1802]*kernel[8];
				ans[1702]<=tmp[1601]*kernel[0]+tmp[1602]*kernel[1]+tmp[1603]*kernel[2]+tmp[1701]*kernel[3]+tmp[1702]*kernel[4]+tmp[1703]*kernel[5]+tmp[1801]*kernel[6]+tmp[1802]*kernel[7]+tmp[1803]*kernel[8];
				ans[1703]<=tmp[1602]*kernel[0]+tmp[1603]*kernel[1]+tmp[1604]*kernel[2]+tmp[1702]*kernel[3]+tmp[1703]*kernel[4]+tmp[1704]*kernel[5]+tmp[1802]*kernel[6]+tmp[1803]*kernel[7]+tmp[1804]*kernel[8];
				ans[1704]<=tmp[1603]*kernel[0]+tmp[1604]*kernel[1]+tmp[1605]*kernel[2]+tmp[1703]*kernel[3]+tmp[1704]*kernel[4]+tmp[1705]*kernel[5]+tmp[1803]*kernel[6]+tmp[1804]*kernel[7]+tmp[1805]*kernel[8];
				ans[1705]<=tmp[1604]*kernel[0]+tmp[1605]*kernel[1]+tmp[1606]*kernel[2]+tmp[1704]*kernel[3]+tmp[1705]*kernel[4]+tmp[1706]*kernel[5]+tmp[1804]*kernel[6]+tmp[1805]*kernel[7]+tmp[1806]*kernel[8];
				ans[1706]<=tmp[1605]*kernel[0]+tmp[1606]*kernel[1]+tmp[1607]*kernel[2]+tmp[1705]*kernel[3]+tmp[1706]*kernel[4]+tmp[1707]*kernel[5]+tmp[1805]*kernel[6]+tmp[1806]*kernel[7]+tmp[1807]*kernel[8];
				ans[1707]<=tmp[1606]*kernel[0]+tmp[1607]*kernel[1]+tmp[1608]*kernel[2]+tmp[1706]*kernel[3]+tmp[1707]*kernel[4]+tmp[1708]*kernel[5]+tmp[1806]*kernel[6]+tmp[1807]*kernel[7]+tmp[1808]*kernel[8];
				ans[1708]<=tmp[1607]*kernel[0]+tmp[1608]*kernel[1]+tmp[1609]*kernel[2]+tmp[1707]*kernel[3]+tmp[1708]*kernel[4]+tmp[1709]*kernel[5]+tmp[1807]*kernel[6]+tmp[1808]*kernel[7]+tmp[1809]*kernel[8];
				ans[1709]<=tmp[1608]*kernel[0]+tmp[1609]*kernel[1]+tmp[1610]*kernel[2]+tmp[1708]*kernel[3]+tmp[1709]*kernel[4]+tmp[1710]*kernel[5]+tmp[1808]*kernel[6]+tmp[1809]*kernel[7]+tmp[1810]*kernel[8];
				ans[1710]<=tmp[1609]*kernel[0]+tmp[1610]*kernel[1]+tmp[1611]*kernel[2]+tmp[1709]*kernel[3]+tmp[1710]*kernel[4]+tmp[1711]*kernel[5]+tmp[1809]*kernel[6]+tmp[1810]*kernel[7]+tmp[1811]*kernel[8];
				ans[1711]<=tmp[1610]*kernel[0]+tmp[1611]*kernel[1]+tmp[1612]*kernel[2]+tmp[1710]*kernel[3]+tmp[1711]*kernel[4]+tmp[1712]*kernel[5]+tmp[1810]*kernel[6]+tmp[1811]*kernel[7]+tmp[1812]*kernel[8];
				ans[1712]<=tmp[1611]*kernel[0]+tmp[1612]*kernel[1]+tmp[1613]*kernel[2]+tmp[1711]*kernel[3]+tmp[1712]*kernel[4]+tmp[1713]*kernel[5]+tmp[1811]*kernel[6]+tmp[1812]*kernel[7]+tmp[1813]*kernel[8];
				ans[1713]<=tmp[1612]*kernel[0]+tmp[1613]*kernel[1]+tmp[1614]*kernel[2]+tmp[1712]*kernel[3]+tmp[1713]*kernel[4]+tmp[1714]*kernel[5]+tmp[1812]*kernel[6]+tmp[1813]*kernel[7]+tmp[1814]*kernel[8];
				ans[1714]<=tmp[1613]*kernel[0]+tmp[1614]*kernel[1]+tmp[1615]*kernel[2]+tmp[1713]*kernel[3]+tmp[1714]*kernel[4]+tmp[1715]*kernel[5]+tmp[1813]*kernel[6]+tmp[1814]*kernel[7]+tmp[1815]*kernel[8];
				ans[1715]<=tmp[1614]*kernel[0]+tmp[1615]*kernel[1]+tmp[1616]*kernel[2]+tmp[1714]*kernel[3]+tmp[1715]*kernel[4]+tmp[1716]*kernel[5]+tmp[1814]*kernel[6]+tmp[1815]*kernel[7]+tmp[1816]*kernel[8];
				ans[1716]<=tmp[1615]*kernel[0]+tmp[1616]*kernel[1]+tmp[1617]*kernel[2]+tmp[1715]*kernel[3]+tmp[1716]*kernel[4]+tmp[1717]*kernel[5]+tmp[1815]*kernel[6]+tmp[1816]*kernel[7]+tmp[1817]*kernel[8];
				ans[1717]<=tmp[1616]*kernel[0]+tmp[1617]*kernel[1]+tmp[1618]*kernel[2]+tmp[1716]*kernel[3]+tmp[1717]*kernel[4]+tmp[1718]*kernel[5]+tmp[1816]*kernel[6]+tmp[1817]*kernel[7]+tmp[1818]*kernel[8];
				ans[1718]<=tmp[1617]*kernel[0]+tmp[1618]*kernel[1]+tmp[1619]*kernel[2]+tmp[1717]*kernel[3]+tmp[1718]*kernel[4]+tmp[1719]*kernel[5]+tmp[1817]*kernel[6]+tmp[1818]*kernel[7]+tmp[1819]*kernel[8];
				ans[1719]<=tmp[1618]*kernel[0]+tmp[1619]*kernel[1]+tmp[1620]*kernel[2]+tmp[1718]*kernel[3]+tmp[1719]*kernel[4]+tmp[1720]*kernel[5]+tmp[1818]*kernel[6]+tmp[1819]*kernel[7]+tmp[1820]*kernel[8];
				ans[1720]<=tmp[1619]*kernel[0]+tmp[1620]*kernel[1]+tmp[1621]*kernel[2]+tmp[1719]*kernel[3]+tmp[1720]*kernel[4]+tmp[1721]*kernel[5]+tmp[1819]*kernel[6]+tmp[1820]*kernel[7]+tmp[1821]*kernel[8];
				ans[1721]<=tmp[1620]*kernel[0]+tmp[1621]*kernel[1]+tmp[1622]*kernel[2]+tmp[1720]*kernel[3]+tmp[1721]*kernel[4]+tmp[1722]*kernel[5]+tmp[1820]*kernel[6]+tmp[1821]*kernel[7]+tmp[1822]*kernel[8];
				ans[1722]<=tmp[1621]*kernel[0]+tmp[1622]*kernel[1]+tmp[1623]*kernel[2]+tmp[1721]*kernel[3]+tmp[1722]*kernel[4]+tmp[1723]*kernel[5]+tmp[1821]*kernel[6]+tmp[1822]*kernel[7]+tmp[1823]*kernel[8];
				ans[1723]<=tmp[1622]*kernel[0]+tmp[1623]*kernel[1]+tmp[1624]*kernel[2]+tmp[1722]*kernel[3]+tmp[1723]*kernel[4]+tmp[1724]*kernel[5]+tmp[1822]*kernel[6]+tmp[1823]*kernel[7]+tmp[1824]*kernel[8];
				ans[1724]<=tmp[1623]*kernel[0]+tmp[1624]*kernel[1]+tmp[1625]*kernel[2]+tmp[1723]*kernel[3]+tmp[1724]*kernel[4]+tmp[1725]*kernel[5]+tmp[1823]*kernel[6]+tmp[1824]*kernel[7]+tmp[1825]*kernel[8];
				ans[1725]<=tmp[1624]*kernel[0]+tmp[1625]*kernel[1]+tmp[1626]*kernel[2]+tmp[1724]*kernel[3]+tmp[1725]*kernel[4]+tmp[1726]*kernel[5]+tmp[1824]*kernel[6]+tmp[1825]*kernel[7]+tmp[1826]*kernel[8];
				ans[1726]<=tmp[1625]*kernel[0]+tmp[1626]*kernel[1]+tmp[1627]*kernel[2]+tmp[1725]*kernel[3]+tmp[1726]*kernel[4]+tmp[1727]*kernel[5]+tmp[1825]*kernel[6]+tmp[1826]*kernel[7]+tmp[1827]*kernel[8];
				ans[1727]<=tmp[1626]*kernel[0]+tmp[1627]*kernel[1]+tmp[1628]*kernel[2]+tmp[1726]*kernel[3]+tmp[1727]*kernel[4]+tmp[1728]*kernel[5]+tmp[1826]*kernel[6]+tmp[1827]*kernel[7]+tmp[1828]*kernel[8];
				ans[1728]<=tmp[1627]*kernel[0]+tmp[1628]*kernel[1]+tmp[1629]*kernel[2]+tmp[1727]*kernel[3]+tmp[1728]*kernel[4]+tmp[1729]*kernel[5]+tmp[1827]*kernel[6]+tmp[1828]*kernel[7]+tmp[1829]*kernel[8];
				ans[1729]<=tmp[1628]*kernel[0]+tmp[1629]*kernel[1]+tmp[1630]*kernel[2]+tmp[1728]*kernel[3]+tmp[1729]*kernel[4]+tmp[1730]*kernel[5]+tmp[1828]*kernel[6]+tmp[1829]*kernel[7]+tmp[1830]*kernel[8];
				ans[1730]<=tmp[1629]*kernel[0]+tmp[1630]*kernel[1]+tmp[1631]*kernel[2]+tmp[1729]*kernel[3]+tmp[1730]*kernel[4]+tmp[1731]*kernel[5]+tmp[1829]*kernel[6]+tmp[1830]*kernel[7]+tmp[1831]*kernel[8];
				ans[1731]<=tmp[1630]*kernel[0]+tmp[1631]*kernel[1]+tmp[1632]*kernel[2]+tmp[1730]*kernel[3]+tmp[1731]*kernel[4]+tmp[1732]*kernel[5]+tmp[1830]*kernel[6]+tmp[1831]*kernel[7]+tmp[1832]*kernel[8];
				ans[1732]<=tmp[1631]*kernel[0]+tmp[1632]*kernel[1]+tmp[1633]*kernel[2]+tmp[1731]*kernel[3]+tmp[1732]*kernel[4]+tmp[1733]*kernel[5]+tmp[1831]*kernel[6]+tmp[1832]*kernel[7]+tmp[1833]*kernel[8];
				ans[1733]<=tmp[1632]*kernel[0]+tmp[1633]*kernel[1]+tmp[1634]*kernel[2]+tmp[1732]*kernel[3]+tmp[1733]*kernel[4]+tmp[1734]*kernel[5]+tmp[1832]*kernel[6]+tmp[1833]*kernel[7]+tmp[1834]*kernel[8];
				ans[1734]<=tmp[1633]*kernel[0]+tmp[1634]*kernel[1]+tmp[1635]*kernel[2]+tmp[1733]*kernel[3]+tmp[1734]*kernel[4]+tmp[1735]*kernel[5]+tmp[1833]*kernel[6]+tmp[1834]*kernel[7]+tmp[1835]*kernel[8];
				ans[1735]<=tmp[1634]*kernel[0]+tmp[1635]*kernel[1]+tmp[1636]*kernel[2]+tmp[1734]*kernel[3]+tmp[1735]*kernel[4]+tmp[1736]*kernel[5]+tmp[1834]*kernel[6]+tmp[1835]*kernel[7]+tmp[1836]*kernel[8];
				ans[1736]<=tmp[1635]*kernel[0]+tmp[1636]*kernel[1]+tmp[1637]*kernel[2]+tmp[1735]*kernel[3]+tmp[1736]*kernel[4]+tmp[1737]*kernel[5]+tmp[1835]*kernel[6]+tmp[1836]*kernel[7]+tmp[1837]*kernel[8];
				ans[1737]<=tmp[1636]*kernel[0]+tmp[1637]*kernel[1]+tmp[1638]*kernel[2]+tmp[1736]*kernel[3]+tmp[1737]*kernel[4]+tmp[1738]*kernel[5]+tmp[1836]*kernel[6]+tmp[1837]*kernel[7]+tmp[1838]*kernel[8];
				ans[1738]<=tmp[1637]*kernel[0]+tmp[1638]*kernel[1]+tmp[1639]*kernel[2]+tmp[1737]*kernel[3]+tmp[1738]*kernel[4]+tmp[1739]*kernel[5]+tmp[1837]*kernel[6]+tmp[1838]*kernel[7]+tmp[1839]*kernel[8];
				ans[1739]<=tmp[1638]*kernel[0]+tmp[1639]*kernel[1]+tmp[1640]*kernel[2]+tmp[1738]*kernel[3]+tmp[1739]*kernel[4]+tmp[1740]*kernel[5]+tmp[1838]*kernel[6]+tmp[1839]*kernel[7]+tmp[1840]*kernel[8];
				ans[1740]<=tmp[1639]*kernel[0]+tmp[1640]*kernel[1]+tmp[1641]*kernel[2]+tmp[1739]*kernel[3]+tmp[1740]*kernel[4]+tmp[1741]*kernel[5]+tmp[1839]*kernel[6]+tmp[1840]*kernel[7]+tmp[1841]*kernel[8];
				ans[1741]<=tmp[1640]*kernel[0]+tmp[1641]*kernel[1]+tmp[1642]*kernel[2]+tmp[1740]*kernel[3]+tmp[1741]*kernel[4]+tmp[1742]*kernel[5]+tmp[1840]*kernel[6]+tmp[1841]*kernel[7]+tmp[1842]*kernel[8];
				ans[1742]<=tmp[1641]*kernel[0]+tmp[1642]*kernel[1]+tmp[1643]*kernel[2]+tmp[1741]*kernel[3]+tmp[1742]*kernel[4]+tmp[1743]*kernel[5]+tmp[1841]*kernel[6]+tmp[1842]*kernel[7]+tmp[1843]*kernel[8];
				ans[1743]<=tmp[1642]*kernel[0]+tmp[1643]*kernel[1]+tmp[1644]*kernel[2]+tmp[1742]*kernel[3]+tmp[1743]*kernel[4]+tmp[1744]*kernel[5]+tmp[1842]*kernel[6]+tmp[1843]*kernel[7]+tmp[1844]*kernel[8];
				ans[1744]<=tmp[1643]*kernel[0]+tmp[1644]*kernel[1]+tmp[1645]*kernel[2]+tmp[1743]*kernel[3]+tmp[1744]*kernel[4]+tmp[1745]*kernel[5]+tmp[1843]*kernel[6]+tmp[1844]*kernel[7]+tmp[1845]*kernel[8];
				ans[1745]<=tmp[1644]*kernel[0]+tmp[1645]*kernel[1]+tmp[1646]*kernel[2]+tmp[1744]*kernel[3]+tmp[1745]*kernel[4]+tmp[1746]*kernel[5]+tmp[1844]*kernel[6]+tmp[1845]*kernel[7]+tmp[1846]*kernel[8];
				ans[1746]<=tmp[1645]*kernel[0]+tmp[1646]*kernel[1]+tmp[1647]*kernel[2]+tmp[1745]*kernel[3]+tmp[1746]*kernel[4]+tmp[1747]*kernel[5]+tmp[1845]*kernel[6]+tmp[1846]*kernel[7]+tmp[1847]*kernel[8];
				ans[1747]<=tmp[1646]*kernel[0]+tmp[1647]*kernel[1]+tmp[1648]*kernel[2]+tmp[1746]*kernel[3]+tmp[1747]*kernel[4]+tmp[1748]*kernel[5]+tmp[1846]*kernel[6]+tmp[1847]*kernel[7]+tmp[1848]*kernel[8];
				ans[1748]<=tmp[1647]*kernel[0]+tmp[1648]*kernel[1]+tmp[1649]*kernel[2]+tmp[1747]*kernel[3]+tmp[1748]*kernel[4]+tmp[1749]*kernel[5]+tmp[1847]*kernel[6]+tmp[1848]*kernel[7]+tmp[1849]*kernel[8];
				ans[1749]<=tmp[1648]*kernel[0]+tmp[1649]*kernel[1]+tmp[1650]*kernel[2]+tmp[1748]*kernel[3]+tmp[1749]*kernel[4]+tmp[1750]*kernel[5]+tmp[1848]*kernel[6]+tmp[1849]*kernel[7]+tmp[1850]*kernel[8];
				ans[1750]<=tmp[1649]*kernel[0]+tmp[1650]*kernel[1]+tmp[1651]*kernel[2]+tmp[1749]*kernel[3]+tmp[1750]*kernel[4]+tmp[1751]*kernel[5]+tmp[1849]*kernel[6]+tmp[1850]*kernel[7]+tmp[1851]*kernel[8];
				ans[1751]<=tmp[1650]*kernel[0]+tmp[1651]*kernel[1]+tmp[1652]*kernel[2]+tmp[1750]*kernel[3]+tmp[1751]*kernel[4]+tmp[1752]*kernel[5]+tmp[1850]*kernel[6]+tmp[1851]*kernel[7]+tmp[1852]*kernel[8];
				ans[1752]<=tmp[1651]*kernel[0]+tmp[1652]*kernel[1]+tmp[1653]*kernel[2]+tmp[1751]*kernel[3]+tmp[1752]*kernel[4]+tmp[1753]*kernel[5]+tmp[1851]*kernel[6]+tmp[1852]*kernel[7]+tmp[1853]*kernel[8];
				ans[1753]<=tmp[1652]*kernel[0]+tmp[1653]*kernel[1]+tmp[1654]*kernel[2]+tmp[1752]*kernel[3]+tmp[1753]*kernel[4]+tmp[1754]*kernel[5]+tmp[1852]*kernel[6]+tmp[1853]*kernel[7]+tmp[1854]*kernel[8];
				ans[1754]<=tmp[1653]*kernel[0]+tmp[1654]*kernel[1]+tmp[1655]*kernel[2]+tmp[1753]*kernel[3]+tmp[1754]*kernel[4]+tmp[1755]*kernel[5]+tmp[1853]*kernel[6]+tmp[1854]*kernel[7]+tmp[1855]*kernel[8];
				ans[1755]<=tmp[1654]*kernel[0]+tmp[1655]*kernel[1]+tmp[1656]*kernel[2]+tmp[1754]*kernel[3]+tmp[1755]*kernel[4]+tmp[1756]*kernel[5]+tmp[1854]*kernel[6]+tmp[1855]*kernel[7]+tmp[1856]*kernel[8];
				ans[1756]<=tmp[1655]*kernel[0]+tmp[1656]*kernel[1]+tmp[1657]*kernel[2]+tmp[1755]*kernel[3]+tmp[1756]*kernel[4]+tmp[1757]*kernel[5]+tmp[1855]*kernel[6]+tmp[1856]*kernel[7]+tmp[1857]*kernel[8];
				ans[1757]<=tmp[1656]*kernel[0]+tmp[1657]*kernel[1]+tmp[1658]*kernel[2]+tmp[1756]*kernel[3]+tmp[1757]*kernel[4]+tmp[1758]*kernel[5]+tmp[1856]*kernel[6]+tmp[1857]*kernel[7]+tmp[1858]*kernel[8];
				ans[1758]<=tmp[1657]*kernel[0]+tmp[1658]*kernel[1]+tmp[1659]*kernel[2]+tmp[1757]*kernel[3]+tmp[1758]*kernel[4]+tmp[1759]*kernel[5]+tmp[1857]*kernel[6]+tmp[1858]*kernel[7]+tmp[1859]*kernel[8];
				ans[1759]<=tmp[1658]*kernel[0]+tmp[1659]*kernel[1]+tmp[1660]*kernel[2]+tmp[1758]*kernel[3]+tmp[1759]*kernel[4]+tmp[1760]*kernel[5]+tmp[1858]*kernel[6]+tmp[1859]*kernel[7]+tmp[1860]*kernel[8];
				ans[1760]<=tmp[1659]*kernel[0]+tmp[1660]*kernel[1]+tmp[1661]*kernel[2]+tmp[1759]*kernel[3]+tmp[1760]*kernel[4]+tmp[1761]*kernel[5]+tmp[1859]*kernel[6]+tmp[1860]*kernel[7]+tmp[1861]*kernel[8];
				ans[1761]<=tmp[1660]*kernel[0]+tmp[1661]*kernel[1]+tmp[1662]*kernel[2]+tmp[1760]*kernel[3]+tmp[1761]*kernel[4]+tmp[1762]*kernel[5]+tmp[1860]*kernel[6]+tmp[1861]*kernel[7]+tmp[1862]*kernel[8];
				ans[1762]<=tmp[1661]*kernel[0]+tmp[1662]*kernel[1]+tmp[1663]*kernel[2]+tmp[1761]*kernel[3]+tmp[1762]*kernel[4]+tmp[1763]*kernel[5]+tmp[1861]*kernel[6]+tmp[1862]*kernel[7]+tmp[1863]*kernel[8];
				ans[1763]<=tmp[1662]*kernel[0]+tmp[1663]*kernel[1]+tmp[1664]*kernel[2]+tmp[1762]*kernel[3]+tmp[1763]*kernel[4]+tmp[1764]*kernel[5]+tmp[1862]*kernel[6]+tmp[1863]*kernel[7]+tmp[1864]*kernel[8];
				ans[1764]<=tmp[1663]*kernel[0]+tmp[1664]*kernel[1]+tmp[1665]*kernel[2]+tmp[1763]*kernel[3]+tmp[1764]*kernel[4]+tmp[1765]*kernel[5]+tmp[1863]*kernel[6]+tmp[1864]*kernel[7]+tmp[1865]*kernel[8];
				ans[1765]<=tmp[1664]*kernel[0]+tmp[1665]*kernel[1]+tmp[1666]*kernel[2]+tmp[1764]*kernel[3]+tmp[1765]*kernel[4]+tmp[1766]*kernel[5]+tmp[1864]*kernel[6]+tmp[1865]*kernel[7]+tmp[1866]*kernel[8];
				ans[1766]<=tmp[1665]*kernel[0]+tmp[1666]*kernel[1]+tmp[1667]*kernel[2]+tmp[1765]*kernel[3]+tmp[1766]*kernel[4]+tmp[1767]*kernel[5]+tmp[1865]*kernel[6]+tmp[1866]*kernel[7]+tmp[1867]*kernel[8];
				ans[1767]<=tmp[1666]*kernel[0]+tmp[1667]*kernel[1]+tmp[1668]*kernel[2]+tmp[1766]*kernel[3]+tmp[1767]*kernel[4]+tmp[1768]*kernel[5]+tmp[1866]*kernel[6]+tmp[1867]*kernel[7]+tmp[1868]*kernel[8];
				ans[1768]<=tmp[1667]*kernel[0]+tmp[1668]*kernel[1]+tmp[1669]*kernel[2]+tmp[1767]*kernel[3]+tmp[1768]*kernel[4]+tmp[1769]*kernel[5]+tmp[1867]*kernel[6]+tmp[1868]*kernel[7]+tmp[1869]*kernel[8];
				ans[1769]<=tmp[1668]*kernel[0]+tmp[1669]*kernel[1]+tmp[1670]*kernel[2]+tmp[1768]*kernel[3]+tmp[1769]*kernel[4]+tmp[1770]*kernel[5]+tmp[1868]*kernel[6]+tmp[1869]*kernel[7]+tmp[1870]*kernel[8];
				ans[1770]<=tmp[1669]*kernel[0]+tmp[1670]*kernel[1]+tmp[1671]*kernel[2]+tmp[1769]*kernel[3]+tmp[1770]*kernel[4]+tmp[1771]*kernel[5]+tmp[1869]*kernel[6]+tmp[1870]*kernel[7]+tmp[1871]*kernel[8];
				ans[1771]<=tmp[1670]*kernel[0]+tmp[1671]*kernel[1]+tmp[1672]*kernel[2]+tmp[1770]*kernel[3]+tmp[1771]*kernel[4]+tmp[1772]*kernel[5]+tmp[1870]*kernel[6]+tmp[1871]*kernel[7]+tmp[1872]*kernel[8];
				ans[1772]<=tmp[1671]*kernel[0]+tmp[1672]*kernel[1]+tmp[1673]*kernel[2]+tmp[1771]*kernel[3]+tmp[1772]*kernel[4]+tmp[1773]*kernel[5]+tmp[1871]*kernel[6]+tmp[1872]*kernel[7]+tmp[1873]*kernel[8];
				ans[1773]<=tmp[1672]*kernel[0]+tmp[1673]*kernel[1]+tmp[1674]*kernel[2]+tmp[1772]*kernel[3]+tmp[1773]*kernel[4]+tmp[1774]*kernel[5]+tmp[1872]*kernel[6]+tmp[1873]*kernel[7]+tmp[1874]*kernel[8];
				ans[1774]<=tmp[1673]*kernel[0]+tmp[1674]*kernel[1]+tmp[1675]*kernel[2]+tmp[1773]*kernel[3]+tmp[1774]*kernel[4]+tmp[1775]*kernel[5]+tmp[1873]*kernel[6]+tmp[1874]*kernel[7]+tmp[1875]*kernel[8];
				ans[1775]<=tmp[1674]*kernel[0]+tmp[1675]*kernel[1]+tmp[1676]*kernel[2]+tmp[1774]*kernel[3]+tmp[1775]*kernel[4]+tmp[1776]*kernel[5]+tmp[1874]*kernel[6]+tmp[1875]*kernel[7]+tmp[1876]*kernel[8];
				ans[1776]<=tmp[1675]*kernel[0]+tmp[1676]*kernel[1]+tmp[1677]*kernel[2]+tmp[1775]*kernel[3]+tmp[1776]*kernel[4]+tmp[1777]*kernel[5]+tmp[1875]*kernel[6]+tmp[1876]*kernel[7]+tmp[1877]*kernel[8];
				ans[1777]<=tmp[1676]*kernel[0]+tmp[1677]*kernel[1]+tmp[1678]*kernel[2]+tmp[1776]*kernel[3]+tmp[1777]*kernel[4]+tmp[1778]*kernel[5]+tmp[1876]*kernel[6]+tmp[1877]*kernel[7]+tmp[1878]*kernel[8];
				ans[1778]<=tmp[1677]*kernel[0]+tmp[1678]*kernel[1]+tmp[1679]*kernel[2]+tmp[1777]*kernel[3]+tmp[1778]*kernel[4]+tmp[1779]*kernel[5]+tmp[1877]*kernel[6]+tmp[1878]*kernel[7]+tmp[1879]*kernel[8];
				ans[1779]<=tmp[1678]*kernel[0]+tmp[1679]*kernel[1]+tmp[1680]*kernel[2]+tmp[1778]*kernel[3]+tmp[1779]*kernel[4]+tmp[1780]*kernel[5]+tmp[1878]*kernel[6]+tmp[1879]*kernel[7]+tmp[1880]*kernel[8];
				ans[1780]<=tmp[1679]*kernel[0]+tmp[1680]*kernel[1]+tmp[1681]*kernel[2]+tmp[1779]*kernel[3]+tmp[1780]*kernel[4]+tmp[1781]*kernel[5]+tmp[1879]*kernel[6]+tmp[1880]*kernel[7]+tmp[1881]*kernel[8];
				ans[1781]<=tmp[1680]*kernel[0]+tmp[1681]*kernel[1]+tmp[1682]*kernel[2]+tmp[1780]*kernel[3]+tmp[1781]*kernel[4]+tmp[1782]*kernel[5]+tmp[1880]*kernel[6]+tmp[1881]*kernel[7]+tmp[1882]*kernel[8];
				ans[1782]<=tmp[1681]*kernel[0]+tmp[1682]*kernel[1]+tmp[1683]*kernel[2]+tmp[1781]*kernel[3]+tmp[1782]*kernel[4]+tmp[1783]*kernel[5]+tmp[1881]*kernel[6]+tmp[1882]*kernel[7]+tmp[1883]*kernel[8];
				ans[1783]<=tmp[1682]*kernel[0]+tmp[1683]*kernel[1]+tmp[1684]*kernel[2]+tmp[1782]*kernel[3]+tmp[1783]*kernel[4]+tmp[1784]*kernel[5]+tmp[1882]*kernel[6]+tmp[1883]*kernel[7]+tmp[1884]*kernel[8];
				ans[1784]<=tmp[1683]*kernel[0]+tmp[1684]*kernel[1]+tmp[1685]*kernel[2]+tmp[1783]*kernel[3]+tmp[1784]*kernel[4]+tmp[1785]*kernel[5]+tmp[1883]*kernel[6]+tmp[1884]*kernel[7]+tmp[1885]*kernel[8];
				ans[1785]<=tmp[1684]*kernel[0]+tmp[1685]*kernel[1]+tmp[1686]*kernel[2]+tmp[1784]*kernel[3]+tmp[1785]*kernel[4]+tmp[1786]*kernel[5]+tmp[1884]*kernel[6]+tmp[1885]*kernel[7]+tmp[1886]*kernel[8];
				ans[1786]<=tmp[1685]*kernel[0]+tmp[1686]*kernel[1]+tmp[1687]*kernel[2]+tmp[1785]*kernel[3]+tmp[1786]*kernel[4]+tmp[1787]*kernel[5]+tmp[1885]*kernel[6]+tmp[1886]*kernel[7]+tmp[1887]*kernel[8];
				ans[1787]<=tmp[1686]*kernel[0]+tmp[1687]*kernel[1]+tmp[1688]*kernel[2]+tmp[1786]*kernel[3]+tmp[1787]*kernel[4]+tmp[1788]*kernel[5]+tmp[1886]*kernel[6]+tmp[1887]*kernel[7]+tmp[1888]*kernel[8];
				ans[1788]<=tmp[1687]*kernel[0]+tmp[1688]*kernel[1]+tmp[1689]*kernel[2]+tmp[1787]*kernel[3]+tmp[1788]*kernel[4]+tmp[1789]*kernel[5]+tmp[1887]*kernel[6]+tmp[1888]*kernel[7]+tmp[1889]*kernel[8];
				ans[1789]<=tmp[1688]*kernel[0]+tmp[1689]*kernel[1]+tmp[1690]*kernel[2]+tmp[1788]*kernel[3]+tmp[1789]*kernel[4]+tmp[1790]*kernel[5]+tmp[1888]*kernel[6]+tmp[1889]*kernel[7]+tmp[1890]*kernel[8];
				ans[1790]<=tmp[1689]*kernel[0]+tmp[1690]*kernel[1]+tmp[1691]*kernel[2]+tmp[1789]*kernel[3]+tmp[1790]*kernel[4]+tmp[1791]*kernel[5]+tmp[1889]*kernel[6]+tmp[1890]*kernel[7]+tmp[1891]*kernel[8];
				ans[1791]<=tmp[1690]*kernel[0]+tmp[1691]*kernel[1]+tmp[1692]*kernel[2]+tmp[1790]*kernel[3]+tmp[1791]*kernel[4]+tmp[1792]*kernel[5]+tmp[1890]*kernel[6]+tmp[1891]*kernel[7]+tmp[1892]*kernel[8];
				ans[1792]<=tmp[1691]*kernel[0]+tmp[1692]*kernel[1]+tmp[1693]*kernel[2]+tmp[1791]*kernel[3]+tmp[1792]*kernel[4]+tmp[1793]*kernel[5]+tmp[1891]*kernel[6]+tmp[1892]*kernel[7]+tmp[1893]*kernel[8];
				ans[1793]<=tmp[1692]*kernel[0]+tmp[1693]*kernel[1]+tmp[1694]*kernel[2]+tmp[1792]*kernel[3]+tmp[1793]*kernel[4]+tmp[1794]*kernel[5]+tmp[1892]*kernel[6]+tmp[1893]*kernel[7]+tmp[1894]*kernel[8];
				ans[1794]<=tmp[1693]*kernel[0]+tmp[1694]*kernel[1]+tmp[1695]*kernel[2]+tmp[1793]*kernel[3]+tmp[1794]*kernel[4]+tmp[1795]*kernel[5]+tmp[1893]*kernel[6]+tmp[1894]*kernel[7]+tmp[1895]*kernel[8];
				ans[1795]<=tmp[1694]*kernel[0]+tmp[1695]*kernel[1]+tmp[1696]*kernel[2]+tmp[1794]*kernel[3]+tmp[1795]*kernel[4]+tmp[1796]*kernel[5]+tmp[1894]*kernel[6]+tmp[1895]*kernel[7]+tmp[1896]*kernel[8];
				ans[1796]<=tmp[1695]*kernel[0]+tmp[1696]*kernel[1]+tmp[1697]*kernel[2]+tmp[1795]*kernel[3]+tmp[1796]*kernel[4]+tmp[1797]*kernel[5]+tmp[1895]*kernel[6]+tmp[1896]*kernel[7]+tmp[1897]*kernel[8];
				ans[1797]<=tmp[1696]*kernel[0]+tmp[1697]*kernel[1]+tmp[1698]*kernel[2]+tmp[1796]*kernel[3]+tmp[1797]*kernel[4]+tmp[1798]*kernel[5]+tmp[1896]*kernel[6]+tmp[1897]*kernel[7]+tmp[1898]*kernel[8];
				ans[1798]<=tmp[1697]*kernel[0]+tmp[1698]*kernel[1]+tmp[1699]*kernel[2]+tmp[1797]*kernel[3]+tmp[1798]*kernel[4]+tmp[1799]*kernel[5]+tmp[1897]*kernel[6]+tmp[1898]*kernel[7]+tmp[1899]*kernel[8];
				ans[1799]<=tmp[1698]*kernel[0]+tmp[1699]*kernel[1]+tmp[1798]*kernel[3]+tmp[1799]*kernel[4]+tmp[1898]*kernel[6]+tmp[1899]*kernel[7];
				ans[1800]<=tmp[1700]*kernel[1]+tmp[1701]*kernel[2]+tmp[1800]*kernel[4]+tmp[1801]*kernel[5]+tmp[1900]*kernel[7]+tmp[1901]*kernel[8];
				ans[1801]<=tmp[1700]*kernel[0]+tmp[1701]*kernel[1]+tmp[1702]*kernel[2]+tmp[1800]*kernel[3]+tmp[1801]*kernel[4]+tmp[1802]*kernel[5]+tmp[1900]*kernel[6]+tmp[1901]*kernel[7]+tmp[1902]*kernel[8];
				ans[1802]<=tmp[1701]*kernel[0]+tmp[1702]*kernel[1]+tmp[1703]*kernel[2]+tmp[1801]*kernel[3]+tmp[1802]*kernel[4]+tmp[1803]*kernel[5]+tmp[1901]*kernel[6]+tmp[1902]*kernel[7]+tmp[1903]*kernel[8];
				ans[1803]<=tmp[1702]*kernel[0]+tmp[1703]*kernel[1]+tmp[1704]*kernel[2]+tmp[1802]*kernel[3]+tmp[1803]*kernel[4]+tmp[1804]*kernel[5]+tmp[1902]*kernel[6]+tmp[1903]*kernel[7]+tmp[1904]*kernel[8];
				ans[1804]<=tmp[1703]*kernel[0]+tmp[1704]*kernel[1]+tmp[1705]*kernel[2]+tmp[1803]*kernel[3]+tmp[1804]*kernel[4]+tmp[1805]*kernel[5]+tmp[1903]*kernel[6]+tmp[1904]*kernel[7]+tmp[1905]*kernel[8];
				ans[1805]<=tmp[1704]*kernel[0]+tmp[1705]*kernel[1]+tmp[1706]*kernel[2]+tmp[1804]*kernel[3]+tmp[1805]*kernel[4]+tmp[1806]*kernel[5]+tmp[1904]*kernel[6]+tmp[1905]*kernel[7]+tmp[1906]*kernel[8];
				ans[1806]<=tmp[1705]*kernel[0]+tmp[1706]*kernel[1]+tmp[1707]*kernel[2]+tmp[1805]*kernel[3]+tmp[1806]*kernel[4]+tmp[1807]*kernel[5]+tmp[1905]*kernel[6]+tmp[1906]*kernel[7]+tmp[1907]*kernel[8];
				ans[1807]<=tmp[1706]*kernel[0]+tmp[1707]*kernel[1]+tmp[1708]*kernel[2]+tmp[1806]*kernel[3]+tmp[1807]*kernel[4]+tmp[1808]*kernel[5]+tmp[1906]*kernel[6]+tmp[1907]*kernel[7]+tmp[1908]*kernel[8];
				ans[1808]<=tmp[1707]*kernel[0]+tmp[1708]*kernel[1]+tmp[1709]*kernel[2]+tmp[1807]*kernel[3]+tmp[1808]*kernel[4]+tmp[1809]*kernel[5]+tmp[1907]*kernel[6]+tmp[1908]*kernel[7]+tmp[1909]*kernel[8];
				ans[1809]<=tmp[1708]*kernel[0]+tmp[1709]*kernel[1]+tmp[1710]*kernel[2]+tmp[1808]*kernel[3]+tmp[1809]*kernel[4]+tmp[1810]*kernel[5]+tmp[1908]*kernel[6]+tmp[1909]*kernel[7]+tmp[1910]*kernel[8];
				ans[1810]<=tmp[1709]*kernel[0]+tmp[1710]*kernel[1]+tmp[1711]*kernel[2]+tmp[1809]*kernel[3]+tmp[1810]*kernel[4]+tmp[1811]*kernel[5]+tmp[1909]*kernel[6]+tmp[1910]*kernel[7]+tmp[1911]*kernel[8];
				ans[1811]<=tmp[1710]*kernel[0]+tmp[1711]*kernel[1]+tmp[1712]*kernel[2]+tmp[1810]*kernel[3]+tmp[1811]*kernel[4]+tmp[1812]*kernel[5]+tmp[1910]*kernel[6]+tmp[1911]*kernel[7]+tmp[1912]*kernel[8];
				ans[1812]<=tmp[1711]*kernel[0]+tmp[1712]*kernel[1]+tmp[1713]*kernel[2]+tmp[1811]*kernel[3]+tmp[1812]*kernel[4]+tmp[1813]*kernel[5]+tmp[1911]*kernel[6]+tmp[1912]*kernel[7]+tmp[1913]*kernel[8];
				ans[1813]<=tmp[1712]*kernel[0]+tmp[1713]*kernel[1]+tmp[1714]*kernel[2]+tmp[1812]*kernel[3]+tmp[1813]*kernel[4]+tmp[1814]*kernel[5]+tmp[1912]*kernel[6]+tmp[1913]*kernel[7]+tmp[1914]*kernel[8];
				ans[1814]<=tmp[1713]*kernel[0]+tmp[1714]*kernel[1]+tmp[1715]*kernel[2]+tmp[1813]*kernel[3]+tmp[1814]*kernel[4]+tmp[1815]*kernel[5]+tmp[1913]*kernel[6]+tmp[1914]*kernel[7]+tmp[1915]*kernel[8];
				ans[1815]<=tmp[1714]*kernel[0]+tmp[1715]*kernel[1]+tmp[1716]*kernel[2]+tmp[1814]*kernel[3]+tmp[1815]*kernel[4]+tmp[1816]*kernel[5]+tmp[1914]*kernel[6]+tmp[1915]*kernel[7]+tmp[1916]*kernel[8];
				ans[1816]<=tmp[1715]*kernel[0]+tmp[1716]*kernel[1]+tmp[1717]*kernel[2]+tmp[1815]*kernel[3]+tmp[1816]*kernel[4]+tmp[1817]*kernel[5]+tmp[1915]*kernel[6]+tmp[1916]*kernel[7]+tmp[1917]*kernel[8];
				ans[1817]<=tmp[1716]*kernel[0]+tmp[1717]*kernel[1]+tmp[1718]*kernel[2]+tmp[1816]*kernel[3]+tmp[1817]*kernel[4]+tmp[1818]*kernel[5]+tmp[1916]*kernel[6]+tmp[1917]*kernel[7]+tmp[1918]*kernel[8];
				ans[1818]<=tmp[1717]*kernel[0]+tmp[1718]*kernel[1]+tmp[1719]*kernel[2]+tmp[1817]*kernel[3]+tmp[1818]*kernel[4]+tmp[1819]*kernel[5]+tmp[1917]*kernel[6]+tmp[1918]*kernel[7]+tmp[1919]*kernel[8];
				ans[1819]<=tmp[1718]*kernel[0]+tmp[1719]*kernel[1]+tmp[1720]*kernel[2]+tmp[1818]*kernel[3]+tmp[1819]*kernel[4]+tmp[1820]*kernel[5]+tmp[1918]*kernel[6]+tmp[1919]*kernel[7]+tmp[1920]*kernel[8];
				ans[1820]<=tmp[1719]*kernel[0]+tmp[1720]*kernel[1]+tmp[1721]*kernel[2]+tmp[1819]*kernel[3]+tmp[1820]*kernel[4]+tmp[1821]*kernel[5]+tmp[1919]*kernel[6]+tmp[1920]*kernel[7]+tmp[1921]*kernel[8];
				ans[1821]<=tmp[1720]*kernel[0]+tmp[1721]*kernel[1]+tmp[1722]*kernel[2]+tmp[1820]*kernel[3]+tmp[1821]*kernel[4]+tmp[1822]*kernel[5]+tmp[1920]*kernel[6]+tmp[1921]*kernel[7]+tmp[1922]*kernel[8];
				ans[1822]<=tmp[1721]*kernel[0]+tmp[1722]*kernel[1]+tmp[1723]*kernel[2]+tmp[1821]*kernel[3]+tmp[1822]*kernel[4]+tmp[1823]*kernel[5]+tmp[1921]*kernel[6]+tmp[1922]*kernel[7]+tmp[1923]*kernel[8];
				ans[1823]<=tmp[1722]*kernel[0]+tmp[1723]*kernel[1]+tmp[1724]*kernel[2]+tmp[1822]*kernel[3]+tmp[1823]*kernel[4]+tmp[1824]*kernel[5]+tmp[1922]*kernel[6]+tmp[1923]*kernel[7]+tmp[1924]*kernel[8];
				ans[1824]<=tmp[1723]*kernel[0]+tmp[1724]*kernel[1]+tmp[1725]*kernel[2]+tmp[1823]*kernel[3]+tmp[1824]*kernel[4]+tmp[1825]*kernel[5]+tmp[1923]*kernel[6]+tmp[1924]*kernel[7]+tmp[1925]*kernel[8];
				ans[1825]<=tmp[1724]*kernel[0]+tmp[1725]*kernel[1]+tmp[1726]*kernel[2]+tmp[1824]*kernel[3]+tmp[1825]*kernel[4]+tmp[1826]*kernel[5]+tmp[1924]*kernel[6]+tmp[1925]*kernel[7]+tmp[1926]*kernel[8];
				ans[1826]<=tmp[1725]*kernel[0]+tmp[1726]*kernel[1]+tmp[1727]*kernel[2]+tmp[1825]*kernel[3]+tmp[1826]*kernel[4]+tmp[1827]*kernel[5]+tmp[1925]*kernel[6]+tmp[1926]*kernel[7]+tmp[1927]*kernel[8];
				ans[1827]<=tmp[1726]*kernel[0]+tmp[1727]*kernel[1]+tmp[1728]*kernel[2]+tmp[1826]*kernel[3]+tmp[1827]*kernel[4]+tmp[1828]*kernel[5]+tmp[1926]*kernel[6]+tmp[1927]*kernel[7]+tmp[1928]*kernel[8];
				ans[1828]<=tmp[1727]*kernel[0]+tmp[1728]*kernel[1]+tmp[1729]*kernel[2]+tmp[1827]*kernel[3]+tmp[1828]*kernel[4]+tmp[1829]*kernel[5]+tmp[1927]*kernel[6]+tmp[1928]*kernel[7]+tmp[1929]*kernel[8];
				ans[1829]<=tmp[1728]*kernel[0]+tmp[1729]*kernel[1]+tmp[1730]*kernel[2]+tmp[1828]*kernel[3]+tmp[1829]*kernel[4]+tmp[1830]*kernel[5]+tmp[1928]*kernel[6]+tmp[1929]*kernel[7]+tmp[1930]*kernel[8];
				ans[1830]<=tmp[1729]*kernel[0]+tmp[1730]*kernel[1]+tmp[1731]*kernel[2]+tmp[1829]*kernel[3]+tmp[1830]*kernel[4]+tmp[1831]*kernel[5]+tmp[1929]*kernel[6]+tmp[1930]*kernel[7]+tmp[1931]*kernel[8];
				ans[1831]<=tmp[1730]*kernel[0]+tmp[1731]*kernel[1]+tmp[1732]*kernel[2]+tmp[1830]*kernel[3]+tmp[1831]*kernel[4]+tmp[1832]*kernel[5]+tmp[1930]*kernel[6]+tmp[1931]*kernel[7]+tmp[1932]*kernel[8];
				ans[1832]<=tmp[1731]*kernel[0]+tmp[1732]*kernel[1]+tmp[1733]*kernel[2]+tmp[1831]*kernel[3]+tmp[1832]*kernel[4]+tmp[1833]*kernel[5]+tmp[1931]*kernel[6]+tmp[1932]*kernel[7]+tmp[1933]*kernel[8];
				ans[1833]<=tmp[1732]*kernel[0]+tmp[1733]*kernel[1]+tmp[1734]*kernel[2]+tmp[1832]*kernel[3]+tmp[1833]*kernel[4]+tmp[1834]*kernel[5]+tmp[1932]*kernel[6]+tmp[1933]*kernel[7]+tmp[1934]*kernel[8];
				ans[1834]<=tmp[1733]*kernel[0]+tmp[1734]*kernel[1]+tmp[1735]*kernel[2]+tmp[1833]*kernel[3]+tmp[1834]*kernel[4]+tmp[1835]*kernel[5]+tmp[1933]*kernel[6]+tmp[1934]*kernel[7]+tmp[1935]*kernel[8];
				ans[1835]<=tmp[1734]*kernel[0]+tmp[1735]*kernel[1]+tmp[1736]*kernel[2]+tmp[1834]*kernel[3]+tmp[1835]*kernel[4]+tmp[1836]*kernel[5]+tmp[1934]*kernel[6]+tmp[1935]*kernel[7]+tmp[1936]*kernel[8];
				ans[1836]<=tmp[1735]*kernel[0]+tmp[1736]*kernel[1]+tmp[1737]*kernel[2]+tmp[1835]*kernel[3]+tmp[1836]*kernel[4]+tmp[1837]*kernel[5]+tmp[1935]*kernel[6]+tmp[1936]*kernel[7]+tmp[1937]*kernel[8];
				ans[1837]<=tmp[1736]*kernel[0]+tmp[1737]*kernel[1]+tmp[1738]*kernel[2]+tmp[1836]*kernel[3]+tmp[1837]*kernel[4]+tmp[1838]*kernel[5]+tmp[1936]*kernel[6]+tmp[1937]*kernel[7]+tmp[1938]*kernel[8];
				ans[1838]<=tmp[1737]*kernel[0]+tmp[1738]*kernel[1]+tmp[1739]*kernel[2]+tmp[1837]*kernel[3]+tmp[1838]*kernel[4]+tmp[1839]*kernel[5]+tmp[1937]*kernel[6]+tmp[1938]*kernel[7]+tmp[1939]*kernel[8];
				ans[1839]<=tmp[1738]*kernel[0]+tmp[1739]*kernel[1]+tmp[1740]*kernel[2]+tmp[1838]*kernel[3]+tmp[1839]*kernel[4]+tmp[1840]*kernel[5]+tmp[1938]*kernel[6]+tmp[1939]*kernel[7]+tmp[1940]*kernel[8];
				ans[1840]<=tmp[1739]*kernel[0]+tmp[1740]*kernel[1]+tmp[1741]*kernel[2]+tmp[1839]*kernel[3]+tmp[1840]*kernel[4]+tmp[1841]*kernel[5]+tmp[1939]*kernel[6]+tmp[1940]*kernel[7]+tmp[1941]*kernel[8];
				ans[1841]<=tmp[1740]*kernel[0]+tmp[1741]*kernel[1]+tmp[1742]*kernel[2]+tmp[1840]*kernel[3]+tmp[1841]*kernel[4]+tmp[1842]*kernel[5]+tmp[1940]*kernel[6]+tmp[1941]*kernel[7]+tmp[1942]*kernel[8];
				ans[1842]<=tmp[1741]*kernel[0]+tmp[1742]*kernel[1]+tmp[1743]*kernel[2]+tmp[1841]*kernel[3]+tmp[1842]*kernel[4]+tmp[1843]*kernel[5]+tmp[1941]*kernel[6]+tmp[1942]*kernel[7]+tmp[1943]*kernel[8];
				ans[1843]<=tmp[1742]*kernel[0]+tmp[1743]*kernel[1]+tmp[1744]*kernel[2]+tmp[1842]*kernel[3]+tmp[1843]*kernel[4]+tmp[1844]*kernel[5]+tmp[1942]*kernel[6]+tmp[1943]*kernel[7]+tmp[1944]*kernel[8];
				ans[1844]<=tmp[1743]*kernel[0]+tmp[1744]*kernel[1]+tmp[1745]*kernel[2]+tmp[1843]*kernel[3]+tmp[1844]*kernel[4]+tmp[1845]*kernel[5]+tmp[1943]*kernel[6]+tmp[1944]*kernel[7]+tmp[1945]*kernel[8];
				ans[1845]<=tmp[1744]*kernel[0]+tmp[1745]*kernel[1]+tmp[1746]*kernel[2]+tmp[1844]*kernel[3]+tmp[1845]*kernel[4]+tmp[1846]*kernel[5]+tmp[1944]*kernel[6]+tmp[1945]*kernel[7]+tmp[1946]*kernel[8];
				ans[1846]<=tmp[1745]*kernel[0]+tmp[1746]*kernel[1]+tmp[1747]*kernel[2]+tmp[1845]*kernel[3]+tmp[1846]*kernel[4]+tmp[1847]*kernel[5]+tmp[1945]*kernel[6]+tmp[1946]*kernel[7]+tmp[1947]*kernel[8];
				ans[1847]<=tmp[1746]*kernel[0]+tmp[1747]*kernel[1]+tmp[1748]*kernel[2]+tmp[1846]*kernel[3]+tmp[1847]*kernel[4]+tmp[1848]*kernel[5]+tmp[1946]*kernel[6]+tmp[1947]*kernel[7]+tmp[1948]*kernel[8];
				ans[1848]<=tmp[1747]*kernel[0]+tmp[1748]*kernel[1]+tmp[1749]*kernel[2]+tmp[1847]*kernel[3]+tmp[1848]*kernel[4]+tmp[1849]*kernel[5]+tmp[1947]*kernel[6]+tmp[1948]*kernel[7]+tmp[1949]*kernel[8];
				ans[1849]<=tmp[1748]*kernel[0]+tmp[1749]*kernel[1]+tmp[1750]*kernel[2]+tmp[1848]*kernel[3]+tmp[1849]*kernel[4]+tmp[1850]*kernel[5]+tmp[1948]*kernel[6]+tmp[1949]*kernel[7]+tmp[1950]*kernel[8];
				ans[1850]<=tmp[1749]*kernel[0]+tmp[1750]*kernel[1]+tmp[1751]*kernel[2]+tmp[1849]*kernel[3]+tmp[1850]*kernel[4]+tmp[1851]*kernel[5]+tmp[1949]*kernel[6]+tmp[1950]*kernel[7]+tmp[1951]*kernel[8];
				ans[1851]<=tmp[1750]*kernel[0]+tmp[1751]*kernel[1]+tmp[1752]*kernel[2]+tmp[1850]*kernel[3]+tmp[1851]*kernel[4]+tmp[1852]*kernel[5]+tmp[1950]*kernel[6]+tmp[1951]*kernel[7]+tmp[1952]*kernel[8];
				ans[1852]<=tmp[1751]*kernel[0]+tmp[1752]*kernel[1]+tmp[1753]*kernel[2]+tmp[1851]*kernel[3]+tmp[1852]*kernel[4]+tmp[1853]*kernel[5]+tmp[1951]*kernel[6]+tmp[1952]*kernel[7]+tmp[1953]*kernel[8];
				ans[1853]<=tmp[1752]*kernel[0]+tmp[1753]*kernel[1]+tmp[1754]*kernel[2]+tmp[1852]*kernel[3]+tmp[1853]*kernel[4]+tmp[1854]*kernel[5]+tmp[1952]*kernel[6]+tmp[1953]*kernel[7]+tmp[1954]*kernel[8];
				ans[1854]<=tmp[1753]*kernel[0]+tmp[1754]*kernel[1]+tmp[1755]*kernel[2]+tmp[1853]*kernel[3]+tmp[1854]*kernel[4]+tmp[1855]*kernel[5]+tmp[1953]*kernel[6]+tmp[1954]*kernel[7]+tmp[1955]*kernel[8];
				ans[1855]<=tmp[1754]*kernel[0]+tmp[1755]*kernel[1]+tmp[1756]*kernel[2]+tmp[1854]*kernel[3]+tmp[1855]*kernel[4]+tmp[1856]*kernel[5]+tmp[1954]*kernel[6]+tmp[1955]*kernel[7]+tmp[1956]*kernel[8];
				ans[1856]<=tmp[1755]*kernel[0]+tmp[1756]*kernel[1]+tmp[1757]*kernel[2]+tmp[1855]*kernel[3]+tmp[1856]*kernel[4]+tmp[1857]*kernel[5]+tmp[1955]*kernel[6]+tmp[1956]*kernel[7]+tmp[1957]*kernel[8];
				ans[1857]<=tmp[1756]*kernel[0]+tmp[1757]*kernel[1]+tmp[1758]*kernel[2]+tmp[1856]*kernel[3]+tmp[1857]*kernel[4]+tmp[1858]*kernel[5]+tmp[1956]*kernel[6]+tmp[1957]*kernel[7]+tmp[1958]*kernel[8];
				ans[1858]<=tmp[1757]*kernel[0]+tmp[1758]*kernel[1]+tmp[1759]*kernel[2]+tmp[1857]*kernel[3]+tmp[1858]*kernel[4]+tmp[1859]*kernel[5]+tmp[1957]*kernel[6]+tmp[1958]*kernel[7]+tmp[1959]*kernel[8];
				ans[1859]<=tmp[1758]*kernel[0]+tmp[1759]*kernel[1]+tmp[1760]*kernel[2]+tmp[1858]*kernel[3]+tmp[1859]*kernel[4]+tmp[1860]*kernel[5]+tmp[1958]*kernel[6]+tmp[1959]*kernel[7]+tmp[1960]*kernel[8];
				ans[1860]<=tmp[1759]*kernel[0]+tmp[1760]*kernel[1]+tmp[1761]*kernel[2]+tmp[1859]*kernel[3]+tmp[1860]*kernel[4]+tmp[1861]*kernel[5]+tmp[1959]*kernel[6]+tmp[1960]*kernel[7]+tmp[1961]*kernel[8];
				ans[1861]<=tmp[1760]*kernel[0]+tmp[1761]*kernel[1]+tmp[1762]*kernel[2]+tmp[1860]*kernel[3]+tmp[1861]*kernel[4]+tmp[1862]*kernel[5]+tmp[1960]*kernel[6]+tmp[1961]*kernel[7]+tmp[1962]*kernel[8];
				ans[1862]<=tmp[1761]*kernel[0]+tmp[1762]*kernel[1]+tmp[1763]*kernel[2]+tmp[1861]*kernel[3]+tmp[1862]*kernel[4]+tmp[1863]*kernel[5]+tmp[1961]*kernel[6]+tmp[1962]*kernel[7]+tmp[1963]*kernel[8];
				ans[1863]<=tmp[1762]*kernel[0]+tmp[1763]*kernel[1]+tmp[1764]*kernel[2]+tmp[1862]*kernel[3]+tmp[1863]*kernel[4]+tmp[1864]*kernel[5]+tmp[1962]*kernel[6]+tmp[1963]*kernel[7]+tmp[1964]*kernel[8];
				ans[1864]<=tmp[1763]*kernel[0]+tmp[1764]*kernel[1]+tmp[1765]*kernel[2]+tmp[1863]*kernel[3]+tmp[1864]*kernel[4]+tmp[1865]*kernel[5]+tmp[1963]*kernel[6]+tmp[1964]*kernel[7]+tmp[1965]*kernel[8];
				ans[1865]<=tmp[1764]*kernel[0]+tmp[1765]*kernel[1]+tmp[1766]*kernel[2]+tmp[1864]*kernel[3]+tmp[1865]*kernel[4]+tmp[1866]*kernel[5]+tmp[1964]*kernel[6]+tmp[1965]*kernel[7]+tmp[1966]*kernel[8];
				ans[1866]<=tmp[1765]*kernel[0]+tmp[1766]*kernel[1]+tmp[1767]*kernel[2]+tmp[1865]*kernel[3]+tmp[1866]*kernel[4]+tmp[1867]*kernel[5]+tmp[1965]*kernel[6]+tmp[1966]*kernel[7]+tmp[1967]*kernel[8];
				ans[1867]<=tmp[1766]*kernel[0]+tmp[1767]*kernel[1]+tmp[1768]*kernel[2]+tmp[1866]*kernel[3]+tmp[1867]*kernel[4]+tmp[1868]*kernel[5]+tmp[1966]*kernel[6]+tmp[1967]*kernel[7]+tmp[1968]*kernel[8];
				ans[1868]<=tmp[1767]*kernel[0]+tmp[1768]*kernel[1]+tmp[1769]*kernel[2]+tmp[1867]*kernel[3]+tmp[1868]*kernel[4]+tmp[1869]*kernel[5]+tmp[1967]*kernel[6]+tmp[1968]*kernel[7]+tmp[1969]*kernel[8];
				ans[1869]<=tmp[1768]*kernel[0]+tmp[1769]*kernel[1]+tmp[1770]*kernel[2]+tmp[1868]*kernel[3]+tmp[1869]*kernel[4]+tmp[1870]*kernel[5]+tmp[1968]*kernel[6]+tmp[1969]*kernel[7]+tmp[1970]*kernel[8];
				ans[1870]<=tmp[1769]*kernel[0]+tmp[1770]*kernel[1]+tmp[1771]*kernel[2]+tmp[1869]*kernel[3]+tmp[1870]*kernel[4]+tmp[1871]*kernel[5]+tmp[1969]*kernel[6]+tmp[1970]*kernel[7]+tmp[1971]*kernel[8];
				ans[1871]<=tmp[1770]*kernel[0]+tmp[1771]*kernel[1]+tmp[1772]*kernel[2]+tmp[1870]*kernel[3]+tmp[1871]*kernel[4]+tmp[1872]*kernel[5]+tmp[1970]*kernel[6]+tmp[1971]*kernel[7]+tmp[1972]*kernel[8];
				ans[1872]<=tmp[1771]*kernel[0]+tmp[1772]*kernel[1]+tmp[1773]*kernel[2]+tmp[1871]*kernel[3]+tmp[1872]*kernel[4]+tmp[1873]*kernel[5]+tmp[1971]*kernel[6]+tmp[1972]*kernel[7]+tmp[1973]*kernel[8];
				ans[1873]<=tmp[1772]*kernel[0]+tmp[1773]*kernel[1]+tmp[1774]*kernel[2]+tmp[1872]*kernel[3]+tmp[1873]*kernel[4]+tmp[1874]*kernel[5]+tmp[1972]*kernel[6]+tmp[1973]*kernel[7]+tmp[1974]*kernel[8];
				ans[1874]<=tmp[1773]*kernel[0]+tmp[1774]*kernel[1]+tmp[1775]*kernel[2]+tmp[1873]*kernel[3]+tmp[1874]*kernel[4]+tmp[1875]*kernel[5]+tmp[1973]*kernel[6]+tmp[1974]*kernel[7]+tmp[1975]*kernel[8];
				ans[1875]<=tmp[1774]*kernel[0]+tmp[1775]*kernel[1]+tmp[1776]*kernel[2]+tmp[1874]*kernel[3]+tmp[1875]*kernel[4]+tmp[1876]*kernel[5]+tmp[1974]*kernel[6]+tmp[1975]*kernel[7]+tmp[1976]*kernel[8];
				ans[1876]<=tmp[1775]*kernel[0]+tmp[1776]*kernel[1]+tmp[1777]*kernel[2]+tmp[1875]*kernel[3]+tmp[1876]*kernel[4]+tmp[1877]*kernel[5]+tmp[1975]*kernel[6]+tmp[1976]*kernel[7]+tmp[1977]*kernel[8];
				ans[1877]<=tmp[1776]*kernel[0]+tmp[1777]*kernel[1]+tmp[1778]*kernel[2]+tmp[1876]*kernel[3]+tmp[1877]*kernel[4]+tmp[1878]*kernel[5]+tmp[1976]*kernel[6]+tmp[1977]*kernel[7]+tmp[1978]*kernel[8];
				ans[1878]<=tmp[1777]*kernel[0]+tmp[1778]*kernel[1]+tmp[1779]*kernel[2]+tmp[1877]*kernel[3]+tmp[1878]*kernel[4]+tmp[1879]*kernel[5]+tmp[1977]*kernel[6]+tmp[1978]*kernel[7]+tmp[1979]*kernel[8];
				ans[1879]<=tmp[1778]*kernel[0]+tmp[1779]*kernel[1]+tmp[1780]*kernel[2]+tmp[1878]*kernel[3]+tmp[1879]*kernel[4]+tmp[1880]*kernel[5]+tmp[1978]*kernel[6]+tmp[1979]*kernel[7]+tmp[1980]*kernel[8];
				ans[1880]<=tmp[1779]*kernel[0]+tmp[1780]*kernel[1]+tmp[1781]*kernel[2]+tmp[1879]*kernel[3]+tmp[1880]*kernel[4]+tmp[1881]*kernel[5]+tmp[1979]*kernel[6]+tmp[1980]*kernel[7]+tmp[1981]*kernel[8];
				ans[1881]<=tmp[1780]*kernel[0]+tmp[1781]*kernel[1]+tmp[1782]*kernel[2]+tmp[1880]*kernel[3]+tmp[1881]*kernel[4]+tmp[1882]*kernel[5]+tmp[1980]*kernel[6]+tmp[1981]*kernel[7]+tmp[1982]*kernel[8];
				ans[1882]<=tmp[1781]*kernel[0]+tmp[1782]*kernel[1]+tmp[1783]*kernel[2]+tmp[1881]*kernel[3]+tmp[1882]*kernel[4]+tmp[1883]*kernel[5]+tmp[1981]*kernel[6]+tmp[1982]*kernel[7]+tmp[1983]*kernel[8];
				ans[1883]<=tmp[1782]*kernel[0]+tmp[1783]*kernel[1]+tmp[1784]*kernel[2]+tmp[1882]*kernel[3]+tmp[1883]*kernel[4]+tmp[1884]*kernel[5]+tmp[1982]*kernel[6]+tmp[1983]*kernel[7]+tmp[1984]*kernel[8];
				ans[1884]<=tmp[1783]*kernel[0]+tmp[1784]*kernel[1]+tmp[1785]*kernel[2]+tmp[1883]*kernel[3]+tmp[1884]*kernel[4]+tmp[1885]*kernel[5]+tmp[1983]*kernel[6]+tmp[1984]*kernel[7]+tmp[1985]*kernel[8];
				ans[1885]<=tmp[1784]*kernel[0]+tmp[1785]*kernel[1]+tmp[1786]*kernel[2]+tmp[1884]*kernel[3]+tmp[1885]*kernel[4]+tmp[1886]*kernel[5]+tmp[1984]*kernel[6]+tmp[1985]*kernel[7]+tmp[1986]*kernel[8];
				ans[1886]<=tmp[1785]*kernel[0]+tmp[1786]*kernel[1]+tmp[1787]*kernel[2]+tmp[1885]*kernel[3]+tmp[1886]*kernel[4]+tmp[1887]*kernel[5]+tmp[1985]*kernel[6]+tmp[1986]*kernel[7]+tmp[1987]*kernel[8];
				ans[1887]<=tmp[1786]*kernel[0]+tmp[1787]*kernel[1]+tmp[1788]*kernel[2]+tmp[1886]*kernel[3]+tmp[1887]*kernel[4]+tmp[1888]*kernel[5]+tmp[1986]*kernel[6]+tmp[1987]*kernel[7]+tmp[1988]*kernel[8];
				ans[1888]<=tmp[1787]*kernel[0]+tmp[1788]*kernel[1]+tmp[1789]*kernel[2]+tmp[1887]*kernel[3]+tmp[1888]*kernel[4]+tmp[1889]*kernel[5]+tmp[1987]*kernel[6]+tmp[1988]*kernel[7]+tmp[1989]*kernel[8];
				ans[1889]<=tmp[1788]*kernel[0]+tmp[1789]*kernel[1]+tmp[1790]*kernel[2]+tmp[1888]*kernel[3]+tmp[1889]*kernel[4]+tmp[1890]*kernel[5]+tmp[1988]*kernel[6]+tmp[1989]*kernel[7]+tmp[1990]*kernel[8];
				ans[1890]<=tmp[1789]*kernel[0]+tmp[1790]*kernel[1]+tmp[1791]*kernel[2]+tmp[1889]*kernel[3]+tmp[1890]*kernel[4]+tmp[1891]*kernel[5]+tmp[1989]*kernel[6]+tmp[1990]*kernel[7]+tmp[1991]*kernel[8];
				ans[1891]<=tmp[1790]*kernel[0]+tmp[1791]*kernel[1]+tmp[1792]*kernel[2]+tmp[1890]*kernel[3]+tmp[1891]*kernel[4]+tmp[1892]*kernel[5]+tmp[1990]*kernel[6]+tmp[1991]*kernel[7]+tmp[1992]*kernel[8];
				ans[1892]<=tmp[1791]*kernel[0]+tmp[1792]*kernel[1]+tmp[1793]*kernel[2]+tmp[1891]*kernel[3]+tmp[1892]*kernel[4]+tmp[1893]*kernel[5]+tmp[1991]*kernel[6]+tmp[1992]*kernel[7]+tmp[1993]*kernel[8];
				ans[1893]<=tmp[1792]*kernel[0]+tmp[1793]*kernel[1]+tmp[1794]*kernel[2]+tmp[1892]*kernel[3]+tmp[1893]*kernel[4]+tmp[1894]*kernel[5]+tmp[1992]*kernel[6]+tmp[1993]*kernel[7]+tmp[1994]*kernel[8];
				ans[1894]<=tmp[1793]*kernel[0]+tmp[1794]*kernel[1]+tmp[1795]*kernel[2]+tmp[1893]*kernel[3]+tmp[1894]*kernel[4]+tmp[1895]*kernel[5]+tmp[1993]*kernel[6]+tmp[1994]*kernel[7]+tmp[1995]*kernel[8];
				ans[1895]<=tmp[1794]*kernel[0]+tmp[1795]*kernel[1]+tmp[1796]*kernel[2]+tmp[1894]*kernel[3]+tmp[1895]*kernel[4]+tmp[1896]*kernel[5]+tmp[1994]*kernel[6]+tmp[1995]*kernel[7]+tmp[1996]*kernel[8];
				ans[1896]<=tmp[1795]*kernel[0]+tmp[1796]*kernel[1]+tmp[1797]*kernel[2]+tmp[1895]*kernel[3]+tmp[1896]*kernel[4]+tmp[1897]*kernel[5]+tmp[1995]*kernel[6]+tmp[1996]*kernel[7]+tmp[1997]*kernel[8];
				ans[1897]<=tmp[1796]*kernel[0]+tmp[1797]*kernel[1]+tmp[1798]*kernel[2]+tmp[1896]*kernel[3]+tmp[1897]*kernel[4]+tmp[1898]*kernel[5]+tmp[1996]*kernel[6]+tmp[1997]*kernel[7]+tmp[1998]*kernel[8];
				ans[1898]<=tmp[1797]*kernel[0]+tmp[1798]*kernel[1]+tmp[1799]*kernel[2]+tmp[1897]*kernel[3]+tmp[1898]*kernel[4]+tmp[1899]*kernel[5]+tmp[1997]*kernel[6]+tmp[1998]*kernel[7]+tmp[1999]*kernel[8];
				ans[1899]<=tmp[1798]*kernel[0]+tmp[1799]*kernel[1]+tmp[1898]*kernel[3]+tmp[1899]*kernel[4]+tmp[1998]*kernel[6]+tmp[1999]*kernel[7];
				ans[1900]<=tmp[1800]*kernel[1]+tmp[1801]*kernel[2]+tmp[1900]*kernel[4]+tmp[1901]*kernel[5]+tmp[2000]*kernel[7]+tmp[2001]*kernel[8];
				ans[1901]<=tmp[1800]*kernel[0]+tmp[1801]*kernel[1]+tmp[1802]*kernel[2]+tmp[1900]*kernel[3]+tmp[1901]*kernel[4]+tmp[1902]*kernel[5]+tmp[2000]*kernel[6]+tmp[2001]*kernel[7]+tmp[2002]*kernel[8];
				ans[1902]<=tmp[1801]*kernel[0]+tmp[1802]*kernel[1]+tmp[1803]*kernel[2]+tmp[1901]*kernel[3]+tmp[1902]*kernel[4]+tmp[1903]*kernel[5]+tmp[2001]*kernel[6]+tmp[2002]*kernel[7]+tmp[2003]*kernel[8];
				ans[1903]<=tmp[1802]*kernel[0]+tmp[1803]*kernel[1]+tmp[1804]*kernel[2]+tmp[1902]*kernel[3]+tmp[1903]*kernel[4]+tmp[1904]*kernel[5]+tmp[2002]*kernel[6]+tmp[2003]*kernel[7]+tmp[2004]*kernel[8];
				ans[1904]<=tmp[1803]*kernel[0]+tmp[1804]*kernel[1]+tmp[1805]*kernel[2]+tmp[1903]*kernel[3]+tmp[1904]*kernel[4]+tmp[1905]*kernel[5]+tmp[2003]*kernel[6]+tmp[2004]*kernel[7]+tmp[2005]*kernel[8];
				ans[1905]<=tmp[1804]*kernel[0]+tmp[1805]*kernel[1]+tmp[1806]*kernel[2]+tmp[1904]*kernel[3]+tmp[1905]*kernel[4]+tmp[1906]*kernel[5]+tmp[2004]*kernel[6]+tmp[2005]*kernel[7]+tmp[2006]*kernel[8];
				ans[1906]<=tmp[1805]*kernel[0]+tmp[1806]*kernel[1]+tmp[1807]*kernel[2]+tmp[1905]*kernel[3]+tmp[1906]*kernel[4]+tmp[1907]*kernel[5]+tmp[2005]*kernel[6]+tmp[2006]*kernel[7]+tmp[2007]*kernel[8];
				ans[1907]<=tmp[1806]*kernel[0]+tmp[1807]*kernel[1]+tmp[1808]*kernel[2]+tmp[1906]*kernel[3]+tmp[1907]*kernel[4]+tmp[1908]*kernel[5]+tmp[2006]*kernel[6]+tmp[2007]*kernel[7]+tmp[2008]*kernel[8];
				ans[1908]<=tmp[1807]*kernel[0]+tmp[1808]*kernel[1]+tmp[1809]*kernel[2]+tmp[1907]*kernel[3]+tmp[1908]*kernel[4]+tmp[1909]*kernel[5]+tmp[2007]*kernel[6]+tmp[2008]*kernel[7]+tmp[2009]*kernel[8];
				ans[1909]<=tmp[1808]*kernel[0]+tmp[1809]*kernel[1]+tmp[1810]*kernel[2]+tmp[1908]*kernel[3]+tmp[1909]*kernel[4]+tmp[1910]*kernel[5]+tmp[2008]*kernel[6]+tmp[2009]*kernel[7]+tmp[2010]*kernel[8];
				ans[1910]<=tmp[1809]*kernel[0]+tmp[1810]*kernel[1]+tmp[1811]*kernel[2]+tmp[1909]*kernel[3]+tmp[1910]*kernel[4]+tmp[1911]*kernel[5]+tmp[2009]*kernel[6]+tmp[2010]*kernel[7]+tmp[2011]*kernel[8];
				ans[1911]<=tmp[1810]*kernel[0]+tmp[1811]*kernel[1]+tmp[1812]*kernel[2]+tmp[1910]*kernel[3]+tmp[1911]*kernel[4]+tmp[1912]*kernel[5]+tmp[2010]*kernel[6]+tmp[2011]*kernel[7]+tmp[2012]*kernel[8];
				ans[1912]<=tmp[1811]*kernel[0]+tmp[1812]*kernel[1]+tmp[1813]*kernel[2]+tmp[1911]*kernel[3]+tmp[1912]*kernel[4]+tmp[1913]*kernel[5]+tmp[2011]*kernel[6]+tmp[2012]*kernel[7]+tmp[2013]*kernel[8];
				ans[1913]<=tmp[1812]*kernel[0]+tmp[1813]*kernel[1]+tmp[1814]*kernel[2]+tmp[1912]*kernel[3]+tmp[1913]*kernel[4]+tmp[1914]*kernel[5]+tmp[2012]*kernel[6]+tmp[2013]*kernel[7]+tmp[2014]*kernel[8];
				ans[1914]<=tmp[1813]*kernel[0]+tmp[1814]*kernel[1]+tmp[1815]*kernel[2]+tmp[1913]*kernel[3]+tmp[1914]*kernel[4]+tmp[1915]*kernel[5]+tmp[2013]*kernel[6]+tmp[2014]*kernel[7]+tmp[2015]*kernel[8];
				ans[1915]<=tmp[1814]*kernel[0]+tmp[1815]*kernel[1]+tmp[1816]*kernel[2]+tmp[1914]*kernel[3]+tmp[1915]*kernel[4]+tmp[1916]*kernel[5]+tmp[2014]*kernel[6]+tmp[2015]*kernel[7]+tmp[2016]*kernel[8];
				ans[1916]<=tmp[1815]*kernel[0]+tmp[1816]*kernel[1]+tmp[1817]*kernel[2]+tmp[1915]*kernel[3]+tmp[1916]*kernel[4]+tmp[1917]*kernel[5]+tmp[2015]*kernel[6]+tmp[2016]*kernel[7]+tmp[2017]*kernel[8];
				ans[1917]<=tmp[1816]*kernel[0]+tmp[1817]*kernel[1]+tmp[1818]*kernel[2]+tmp[1916]*kernel[3]+tmp[1917]*kernel[4]+tmp[1918]*kernel[5]+tmp[2016]*kernel[6]+tmp[2017]*kernel[7]+tmp[2018]*kernel[8];
				ans[1918]<=tmp[1817]*kernel[0]+tmp[1818]*kernel[1]+tmp[1819]*kernel[2]+tmp[1917]*kernel[3]+tmp[1918]*kernel[4]+tmp[1919]*kernel[5]+tmp[2017]*kernel[6]+tmp[2018]*kernel[7]+tmp[2019]*kernel[8];
				ans[1919]<=tmp[1818]*kernel[0]+tmp[1819]*kernel[1]+tmp[1820]*kernel[2]+tmp[1918]*kernel[3]+tmp[1919]*kernel[4]+tmp[1920]*kernel[5]+tmp[2018]*kernel[6]+tmp[2019]*kernel[7]+tmp[2020]*kernel[8];
				ans[1920]<=tmp[1819]*kernel[0]+tmp[1820]*kernel[1]+tmp[1821]*kernel[2]+tmp[1919]*kernel[3]+tmp[1920]*kernel[4]+tmp[1921]*kernel[5]+tmp[2019]*kernel[6]+tmp[2020]*kernel[7]+tmp[2021]*kernel[8];
				ans[1921]<=tmp[1820]*kernel[0]+tmp[1821]*kernel[1]+tmp[1822]*kernel[2]+tmp[1920]*kernel[3]+tmp[1921]*kernel[4]+tmp[1922]*kernel[5]+tmp[2020]*kernel[6]+tmp[2021]*kernel[7]+tmp[2022]*kernel[8];
				ans[1922]<=tmp[1821]*kernel[0]+tmp[1822]*kernel[1]+tmp[1823]*kernel[2]+tmp[1921]*kernel[3]+tmp[1922]*kernel[4]+tmp[1923]*kernel[5]+tmp[2021]*kernel[6]+tmp[2022]*kernel[7]+tmp[2023]*kernel[8];
				ans[1923]<=tmp[1822]*kernel[0]+tmp[1823]*kernel[1]+tmp[1824]*kernel[2]+tmp[1922]*kernel[3]+tmp[1923]*kernel[4]+tmp[1924]*kernel[5]+tmp[2022]*kernel[6]+tmp[2023]*kernel[7]+tmp[2024]*kernel[8];
				ans[1924]<=tmp[1823]*kernel[0]+tmp[1824]*kernel[1]+tmp[1825]*kernel[2]+tmp[1923]*kernel[3]+tmp[1924]*kernel[4]+tmp[1925]*kernel[5]+tmp[2023]*kernel[6]+tmp[2024]*kernel[7]+tmp[2025]*kernel[8];
				ans[1925]<=tmp[1824]*kernel[0]+tmp[1825]*kernel[1]+tmp[1826]*kernel[2]+tmp[1924]*kernel[3]+tmp[1925]*kernel[4]+tmp[1926]*kernel[5]+tmp[2024]*kernel[6]+tmp[2025]*kernel[7]+tmp[2026]*kernel[8];
				ans[1926]<=tmp[1825]*kernel[0]+tmp[1826]*kernel[1]+tmp[1827]*kernel[2]+tmp[1925]*kernel[3]+tmp[1926]*kernel[4]+tmp[1927]*kernel[5]+tmp[2025]*kernel[6]+tmp[2026]*kernel[7]+tmp[2027]*kernel[8];
				ans[1927]<=tmp[1826]*kernel[0]+tmp[1827]*kernel[1]+tmp[1828]*kernel[2]+tmp[1926]*kernel[3]+tmp[1927]*kernel[4]+tmp[1928]*kernel[5]+tmp[2026]*kernel[6]+tmp[2027]*kernel[7]+tmp[2028]*kernel[8];
				ans[1928]<=tmp[1827]*kernel[0]+tmp[1828]*kernel[1]+tmp[1829]*kernel[2]+tmp[1927]*kernel[3]+tmp[1928]*kernel[4]+tmp[1929]*kernel[5]+tmp[2027]*kernel[6]+tmp[2028]*kernel[7]+tmp[2029]*kernel[8];
				ans[1929]<=tmp[1828]*kernel[0]+tmp[1829]*kernel[1]+tmp[1830]*kernel[2]+tmp[1928]*kernel[3]+tmp[1929]*kernel[4]+tmp[1930]*kernel[5]+tmp[2028]*kernel[6]+tmp[2029]*kernel[7]+tmp[2030]*kernel[8];
				ans[1930]<=tmp[1829]*kernel[0]+tmp[1830]*kernel[1]+tmp[1831]*kernel[2]+tmp[1929]*kernel[3]+tmp[1930]*kernel[4]+tmp[1931]*kernel[5]+tmp[2029]*kernel[6]+tmp[2030]*kernel[7]+tmp[2031]*kernel[8];
				ans[1931]<=tmp[1830]*kernel[0]+tmp[1831]*kernel[1]+tmp[1832]*kernel[2]+tmp[1930]*kernel[3]+tmp[1931]*kernel[4]+tmp[1932]*kernel[5]+tmp[2030]*kernel[6]+tmp[2031]*kernel[7]+tmp[2032]*kernel[8];
				ans[1932]<=tmp[1831]*kernel[0]+tmp[1832]*kernel[1]+tmp[1833]*kernel[2]+tmp[1931]*kernel[3]+tmp[1932]*kernel[4]+tmp[1933]*kernel[5]+tmp[2031]*kernel[6]+tmp[2032]*kernel[7]+tmp[2033]*kernel[8];
				ans[1933]<=tmp[1832]*kernel[0]+tmp[1833]*kernel[1]+tmp[1834]*kernel[2]+tmp[1932]*kernel[3]+tmp[1933]*kernel[4]+tmp[1934]*kernel[5]+tmp[2032]*kernel[6]+tmp[2033]*kernel[7]+tmp[2034]*kernel[8];
				ans[1934]<=tmp[1833]*kernel[0]+tmp[1834]*kernel[1]+tmp[1835]*kernel[2]+tmp[1933]*kernel[3]+tmp[1934]*kernel[4]+tmp[1935]*kernel[5]+tmp[2033]*kernel[6]+tmp[2034]*kernel[7]+tmp[2035]*kernel[8];
				ans[1935]<=tmp[1834]*kernel[0]+tmp[1835]*kernel[1]+tmp[1836]*kernel[2]+tmp[1934]*kernel[3]+tmp[1935]*kernel[4]+tmp[1936]*kernel[5]+tmp[2034]*kernel[6]+tmp[2035]*kernel[7]+tmp[2036]*kernel[8];
				ans[1936]<=tmp[1835]*kernel[0]+tmp[1836]*kernel[1]+tmp[1837]*kernel[2]+tmp[1935]*kernel[3]+tmp[1936]*kernel[4]+tmp[1937]*kernel[5]+tmp[2035]*kernel[6]+tmp[2036]*kernel[7]+tmp[2037]*kernel[8];
				ans[1937]<=tmp[1836]*kernel[0]+tmp[1837]*kernel[1]+tmp[1838]*kernel[2]+tmp[1936]*kernel[3]+tmp[1937]*kernel[4]+tmp[1938]*kernel[5]+tmp[2036]*kernel[6]+tmp[2037]*kernel[7]+tmp[2038]*kernel[8];
				ans[1938]<=tmp[1837]*kernel[0]+tmp[1838]*kernel[1]+tmp[1839]*kernel[2]+tmp[1937]*kernel[3]+tmp[1938]*kernel[4]+tmp[1939]*kernel[5]+tmp[2037]*kernel[6]+tmp[2038]*kernel[7]+tmp[2039]*kernel[8];
				ans[1939]<=tmp[1838]*kernel[0]+tmp[1839]*kernel[1]+tmp[1840]*kernel[2]+tmp[1938]*kernel[3]+tmp[1939]*kernel[4]+tmp[1940]*kernel[5]+tmp[2038]*kernel[6]+tmp[2039]*kernel[7]+tmp[2040]*kernel[8];
				ans[1940]<=tmp[1839]*kernel[0]+tmp[1840]*kernel[1]+tmp[1841]*kernel[2]+tmp[1939]*kernel[3]+tmp[1940]*kernel[4]+tmp[1941]*kernel[5]+tmp[2039]*kernel[6]+tmp[2040]*kernel[7]+tmp[2041]*kernel[8];
				ans[1941]<=tmp[1840]*kernel[0]+tmp[1841]*kernel[1]+tmp[1842]*kernel[2]+tmp[1940]*kernel[3]+tmp[1941]*kernel[4]+tmp[1942]*kernel[5]+tmp[2040]*kernel[6]+tmp[2041]*kernel[7]+tmp[2042]*kernel[8];
				ans[1942]<=tmp[1841]*kernel[0]+tmp[1842]*kernel[1]+tmp[1843]*kernel[2]+tmp[1941]*kernel[3]+tmp[1942]*kernel[4]+tmp[1943]*kernel[5]+tmp[2041]*kernel[6]+tmp[2042]*kernel[7]+tmp[2043]*kernel[8];
				ans[1943]<=tmp[1842]*kernel[0]+tmp[1843]*kernel[1]+tmp[1844]*kernel[2]+tmp[1942]*kernel[3]+tmp[1943]*kernel[4]+tmp[1944]*kernel[5]+tmp[2042]*kernel[6]+tmp[2043]*kernel[7]+tmp[2044]*kernel[8];
				ans[1944]<=tmp[1843]*kernel[0]+tmp[1844]*kernel[1]+tmp[1845]*kernel[2]+tmp[1943]*kernel[3]+tmp[1944]*kernel[4]+tmp[1945]*kernel[5]+tmp[2043]*kernel[6]+tmp[2044]*kernel[7]+tmp[2045]*kernel[8];
				ans[1945]<=tmp[1844]*kernel[0]+tmp[1845]*kernel[1]+tmp[1846]*kernel[2]+tmp[1944]*kernel[3]+tmp[1945]*kernel[4]+tmp[1946]*kernel[5]+tmp[2044]*kernel[6]+tmp[2045]*kernel[7]+tmp[2046]*kernel[8];
				ans[1946]<=tmp[1845]*kernel[0]+tmp[1846]*kernel[1]+tmp[1847]*kernel[2]+tmp[1945]*kernel[3]+tmp[1946]*kernel[4]+tmp[1947]*kernel[5]+tmp[2045]*kernel[6]+tmp[2046]*kernel[7]+tmp[2047]*kernel[8];
				ans[1947]<=tmp[1846]*kernel[0]+tmp[1847]*kernel[1]+tmp[1848]*kernel[2]+tmp[1946]*kernel[3]+tmp[1947]*kernel[4]+tmp[1948]*kernel[5]+tmp[2046]*kernel[6]+tmp[2047]*kernel[7]+tmp[2048]*kernel[8];
				ans[1948]<=tmp[1847]*kernel[0]+tmp[1848]*kernel[1]+tmp[1849]*kernel[2]+tmp[1947]*kernel[3]+tmp[1948]*kernel[4]+tmp[1949]*kernel[5]+tmp[2047]*kernel[6]+tmp[2048]*kernel[7]+tmp[2049]*kernel[8];
				ans[1949]<=tmp[1848]*kernel[0]+tmp[1849]*kernel[1]+tmp[1850]*kernel[2]+tmp[1948]*kernel[3]+tmp[1949]*kernel[4]+tmp[1950]*kernel[5]+tmp[2048]*kernel[6]+tmp[2049]*kernel[7]+tmp[2050]*kernel[8];
				ans[1950]<=tmp[1849]*kernel[0]+tmp[1850]*kernel[1]+tmp[1851]*kernel[2]+tmp[1949]*kernel[3]+tmp[1950]*kernel[4]+tmp[1951]*kernel[5]+tmp[2049]*kernel[6]+tmp[2050]*kernel[7]+tmp[2051]*kernel[8];
				ans[1951]<=tmp[1850]*kernel[0]+tmp[1851]*kernel[1]+tmp[1852]*kernel[2]+tmp[1950]*kernel[3]+tmp[1951]*kernel[4]+tmp[1952]*kernel[5]+tmp[2050]*kernel[6]+tmp[2051]*kernel[7]+tmp[2052]*kernel[8];
				ans[1952]<=tmp[1851]*kernel[0]+tmp[1852]*kernel[1]+tmp[1853]*kernel[2]+tmp[1951]*kernel[3]+tmp[1952]*kernel[4]+tmp[1953]*kernel[5]+tmp[2051]*kernel[6]+tmp[2052]*kernel[7]+tmp[2053]*kernel[8];
				ans[1953]<=tmp[1852]*kernel[0]+tmp[1853]*kernel[1]+tmp[1854]*kernel[2]+tmp[1952]*kernel[3]+tmp[1953]*kernel[4]+tmp[1954]*kernel[5]+tmp[2052]*kernel[6]+tmp[2053]*kernel[7]+tmp[2054]*kernel[8];
				ans[1954]<=tmp[1853]*kernel[0]+tmp[1854]*kernel[1]+tmp[1855]*kernel[2]+tmp[1953]*kernel[3]+tmp[1954]*kernel[4]+tmp[1955]*kernel[5]+tmp[2053]*kernel[6]+tmp[2054]*kernel[7]+tmp[2055]*kernel[8];
				ans[1955]<=tmp[1854]*kernel[0]+tmp[1855]*kernel[1]+tmp[1856]*kernel[2]+tmp[1954]*kernel[3]+tmp[1955]*kernel[4]+tmp[1956]*kernel[5]+tmp[2054]*kernel[6]+tmp[2055]*kernel[7]+tmp[2056]*kernel[8];
				ans[1956]<=tmp[1855]*kernel[0]+tmp[1856]*kernel[1]+tmp[1857]*kernel[2]+tmp[1955]*kernel[3]+tmp[1956]*kernel[4]+tmp[1957]*kernel[5]+tmp[2055]*kernel[6]+tmp[2056]*kernel[7]+tmp[2057]*kernel[8];
				ans[1957]<=tmp[1856]*kernel[0]+tmp[1857]*kernel[1]+tmp[1858]*kernel[2]+tmp[1956]*kernel[3]+tmp[1957]*kernel[4]+tmp[1958]*kernel[5]+tmp[2056]*kernel[6]+tmp[2057]*kernel[7]+tmp[2058]*kernel[8];
				ans[1958]<=tmp[1857]*kernel[0]+tmp[1858]*kernel[1]+tmp[1859]*kernel[2]+tmp[1957]*kernel[3]+tmp[1958]*kernel[4]+tmp[1959]*kernel[5]+tmp[2057]*kernel[6]+tmp[2058]*kernel[7]+tmp[2059]*kernel[8];
				ans[1959]<=tmp[1858]*kernel[0]+tmp[1859]*kernel[1]+tmp[1860]*kernel[2]+tmp[1958]*kernel[3]+tmp[1959]*kernel[4]+tmp[1960]*kernel[5]+tmp[2058]*kernel[6]+tmp[2059]*kernel[7]+tmp[2060]*kernel[8];
				ans[1960]<=tmp[1859]*kernel[0]+tmp[1860]*kernel[1]+tmp[1861]*kernel[2]+tmp[1959]*kernel[3]+tmp[1960]*kernel[4]+tmp[1961]*kernel[5]+tmp[2059]*kernel[6]+tmp[2060]*kernel[7]+tmp[2061]*kernel[8];
				ans[1961]<=tmp[1860]*kernel[0]+tmp[1861]*kernel[1]+tmp[1862]*kernel[2]+tmp[1960]*kernel[3]+tmp[1961]*kernel[4]+tmp[1962]*kernel[5]+tmp[2060]*kernel[6]+tmp[2061]*kernel[7]+tmp[2062]*kernel[8];
				ans[1962]<=tmp[1861]*kernel[0]+tmp[1862]*kernel[1]+tmp[1863]*kernel[2]+tmp[1961]*kernel[3]+tmp[1962]*kernel[4]+tmp[1963]*kernel[5]+tmp[2061]*kernel[6]+tmp[2062]*kernel[7]+tmp[2063]*kernel[8];
				ans[1963]<=tmp[1862]*kernel[0]+tmp[1863]*kernel[1]+tmp[1864]*kernel[2]+tmp[1962]*kernel[3]+tmp[1963]*kernel[4]+tmp[1964]*kernel[5]+tmp[2062]*kernel[6]+tmp[2063]*kernel[7]+tmp[2064]*kernel[8];
				ans[1964]<=tmp[1863]*kernel[0]+tmp[1864]*kernel[1]+tmp[1865]*kernel[2]+tmp[1963]*kernel[3]+tmp[1964]*kernel[4]+tmp[1965]*kernel[5]+tmp[2063]*kernel[6]+tmp[2064]*kernel[7]+tmp[2065]*kernel[8];
				ans[1965]<=tmp[1864]*kernel[0]+tmp[1865]*kernel[1]+tmp[1866]*kernel[2]+tmp[1964]*kernel[3]+tmp[1965]*kernel[4]+tmp[1966]*kernel[5]+tmp[2064]*kernel[6]+tmp[2065]*kernel[7]+tmp[2066]*kernel[8];
				ans[1966]<=tmp[1865]*kernel[0]+tmp[1866]*kernel[1]+tmp[1867]*kernel[2]+tmp[1965]*kernel[3]+tmp[1966]*kernel[4]+tmp[1967]*kernel[5]+tmp[2065]*kernel[6]+tmp[2066]*kernel[7]+tmp[2067]*kernel[8];
				ans[1967]<=tmp[1866]*kernel[0]+tmp[1867]*kernel[1]+tmp[1868]*kernel[2]+tmp[1966]*kernel[3]+tmp[1967]*kernel[4]+tmp[1968]*kernel[5]+tmp[2066]*kernel[6]+tmp[2067]*kernel[7]+tmp[2068]*kernel[8];
				ans[1968]<=tmp[1867]*kernel[0]+tmp[1868]*kernel[1]+tmp[1869]*kernel[2]+tmp[1967]*kernel[3]+tmp[1968]*kernel[4]+tmp[1969]*kernel[5]+tmp[2067]*kernel[6]+tmp[2068]*kernel[7]+tmp[2069]*kernel[8];
				ans[1969]<=tmp[1868]*kernel[0]+tmp[1869]*kernel[1]+tmp[1870]*kernel[2]+tmp[1968]*kernel[3]+tmp[1969]*kernel[4]+tmp[1970]*kernel[5]+tmp[2068]*kernel[6]+tmp[2069]*kernel[7]+tmp[2070]*kernel[8];
				ans[1970]<=tmp[1869]*kernel[0]+tmp[1870]*kernel[1]+tmp[1871]*kernel[2]+tmp[1969]*kernel[3]+tmp[1970]*kernel[4]+tmp[1971]*kernel[5]+tmp[2069]*kernel[6]+tmp[2070]*kernel[7]+tmp[2071]*kernel[8];
				ans[1971]<=tmp[1870]*kernel[0]+tmp[1871]*kernel[1]+tmp[1872]*kernel[2]+tmp[1970]*kernel[3]+tmp[1971]*kernel[4]+tmp[1972]*kernel[5]+tmp[2070]*kernel[6]+tmp[2071]*kernel[7]+tmp[2072]*kernel[8];
				ans[1972]<=tmp[1871]*kernel[0]+tmp[1872]*kernel[1]+tmp[1873]*kernel[2]+tmp[1971]*kernel[3]+tmp[1972]*kernel[4]+tmp[1973]*kernel[5]+tmp[2071]*kernel[6]+tmp[2072]*kernel[7]+tmp[2073]*kernel[8];
				ans[1973]<=tmp[1872]*kernel[0]+tmp[1873]*kernel[1]+tmp[1874]*kernel[2]+tmp[1972]*kernel[3]+tmp[1973]*kernel[4]+tmp[1974]*kernel[5]+tmp[2072]*kernel[6]+tmp[2073]*kernel[7]+tmp[2074]*kernel[8];
				ans[1974]<=tmp[1873]*kernel[0]+tmp[1874]*kernel[1]+tmp[1875]*kernel[2]+tmp[1973]*kernel[3]+tmp[1974]*kernel[4]+tmp[1975]*kernel[5]+tmp[2073]*kernel[6]+tmp[2074]*kernel[7]+tmp[2075]*kernel[8];
				ans[1975]<=tmp[1874]*kernel[0]+tmp[1875]*kernel[1]+tmp[1876]*kernel[2]+tmp[1974]*kernel[3]+tmp[1975]*kernel[4]+tmp[1976]*kernel[5]+tmp[2074]*kernel[6]+tmp[2075]*kernel[7]+tmp[2076]*kernel[8];
				ans[1976]<=tmp[1875]*kernel[0]+tmp[1876]*kernel[1]+tmp[1877]*kernel[2]+tmp[1975]*kernel[3]+tmp[1976]*kernel[4]+tmp[1977]*kernel[5]+tmp[2075]*kernel[6]+tmp[2076]*kernel[7]+tmp[2077]*kernel[8];
				ans[1977]<=tmp[1876]*kernel[0]+tmp[1877]*kernel[1]+tmp[1878]*kernel[2]+tmp[1976]*kernel[3]+tmp[1977]*kernel[4]+tmp[1978]*kernel[5]+tmp[2076]*kernel[6]+tmp[2077]*kernel[7]+tmp[2078]*kernel[8];
				ans[1978]<=tmp[1877]*kernel[0]+tmp[1878]*kernel[1]+tmp[1879]*kernel[2]+tmp[1977]*kernel[3]+tmp[1978]*kernel[4]+tmp[1979]*kernel[5]+tmp[2077]*kernel[6]+tmp[2078]*kernel[7]+tmp[2079]*kernel[8];
				ans[1979]<=tmp[1878]*kernel[0]+tmp[1879]*kernel[1]+tmp[1880]*kernel[2]+tmp[1978]*kernel[3]+tmp[1979]*kernel[4]+tmp[1980]*kernel[5]+tmp[2078]*kernel[6]+tmp[2079]*kernel[7]+tmp[2080]*kernel[8];
				ans[1980]<=tmp[1879]*kernel[0]+tmp[1880]*kernel[1]+tmp[1881]*kernel[2]+tmp[1979]*kernel[3]+tmp[1980]*kernel[4]+tmp[1981]*kernel[5]+tmp[2079]*kernel[6]+tmp[2080]*kernel[7]+tmp[2081]*kernel[8];
				ans[1981]<=tmp[1880]*kernel[0]+tmp[1881]*kernel[1]+tmp[1882]*kernel[2]+tmp[1980]*kernel[3]+tmp[1981]*kernel[4]+tmp[1982]*kernel[5]+tmp[2080]*kernel[6]+tmp[2081]*kernel[7]+tmp[2082]*kernel[8];
				ans[1982]<=tmp[1881]*kernel[0]+tmp[1882]*kernel[1]+tmp[1883]*kernel[2]+tmp[1981]*kernel[3]+tmp[1982]*kernel[4]+tmp[1983]*kernel[5]+tmp[2081]*kernel[6]+tmp[2082]*kernel[7]+tmp[2083]*kernel[8];
				ans[1983]<=tmp[1882]*kernel[0]+tmp[1883]*kernel[1]+tmp[1884]*kernel[2]+tmp[1982]*kernel[3]+tmp[1983]*kernel[4]+tmp[1984]*kernel[5]+tmp[2082]*kernel[6]+tmp[2083]*kernel[7]+tmp[2084]*kernel[8];
				ans[1984]<=tmp[1883]*kernel[0]+tmp[1884]*kernel[1]+tmp[1885]*kernel[2]+tmp[1983]*kernel[3]+tmp[1984]*kernel[4]+tmp[1985]*kernel[5]+tmp[2083]*kernel[6]+tmp[2084]*kernel[7]+tmp[2085]*kernel[8];
				ans[1985]<=tmp[1884]*kernel[0]+tmp[1885]*kernel[1]+tmp[1886]*kernel[2]+tmp[1984]*kernel[3]+tmp[1985]*kernel[4]+tmp[1986]*kernel[5]+tmp[2084]*kernel[6]+tmp[2085]*kernel[7]+tmp[2086]*kernel[8];
				ans[1986]<=tmp[1885]*kernel[0]+tmp[1886]*kernel[1]+tmp[1887]*kernel[2]+tmp[1985]*kernel[3]+tmp[1986]*kernel[4]+tmp[1987]*kernel[5]+tmp[2085]*kernel[6]+tmp[2086]*kernel[7]+tmp[2087]*kernel[8];
				ans[1987]<=tmp[1886]*kernel[0]+tmp[1887]*kernel[1]+tmp[1888]*kernel[2]+tmp[1986]*kernel[3]+tmp[1987]*kernel[4]+tmp[1988]*kernel[5]+tmp[2086]*kernel[6]+tmp[2087]*kernel[7]+tmp[2088]*kernel[8];
				ans[1988]<=tmp[1887]*kernel[0]+tmp[1888]*kernel[1]+tmp[1889]*kernel[2]+tmp[1987]*kernel[3]+tmp[1988]*kernel[4]+tmp[1989]*kernel[5]+tmp[2087]*kernel[6]+tmp[2088]*kernel[7]+tmp[2089]*kernel[8];
				ans[1989]<=tmp[1888]*kernel[0]+tmp[1889]*kernel[1]+tmp[1890]*kernel[2]+tmp[1988]*kernel[3]+tmp[1989]*kernel[4]+tmp[1990]*kernel[5]+tmp[2088]*kernel[6]+tmp[2089]*kernel[7]+tmp[2090]*kernel[8];
				ans[1990]<=tmp[1889]*kernel[0]+tmp[1890]*kernel[1]+tmp[1891]*kernel[2]+tmp[1989]*kernel[3]+tmp[1990]*kernel[4]+tmp[1991]*kernel[5]+tmp[2089]*kernel[6]+tmp[2090]*kernel[7]+tmp[2091]*kernel[8];
				ans[1991]<=tmp[1890]*kernel[0]+tmp[1891]*kernel[1]+tmp[1892]*kernel[2]+tmp[1990]*kernel[3]+tmp[1991]*kernel[4]+tmp[1992]*kernel[5]+tmp[2090]*kernel[6]+tmp[2091]*kernel[7]+tmp[2092]*kernel[8];
				ans[1992]<=tmp[1891]*kernel[0]+tmp[1892]*kernel[1]+tmp[1893]*kernel[2]+tmp[1991]*kernel[3]+tmp[1992]*kernel[4]+tmp[1993]*kernel[5]+tmp[2091]*kernel[6]+tmp[2092]*kernel[7]+tmp[2093]*kernel[8];
				ans[1993]<=tmp[1892]*kernel[0]+tmp[1893]*kernel[1]+tmp[1894]*kernel[2]+tmp[1992]*kernel[3]+tmp[1993]*kernel[4]+tmp[1994]*kernel[5]+tmp[2092]*kernel[6]+tmp[2093]*kernel[7]+tmp[2094]*kernel[8];
				ans[1994]<=tmp[1893]*kernel[0]+tmp[1894]*kernel[1]+tmp[1895]*kernel[2]+tmp[1993]*kernel[3]+tmp[1994]*kernel[4]+tmp[1995]*kernel[5]+tmp[2093]*kernel[6]+tmp[2094]*kernel[7]+tmp[2095]*kernel[8];
				ans[1995]<=tmp[1894]*kernel[0]+tmp[1895]*kernel[1]+tmp[1896]*kernel[2]+tmp[1994]*kernel[3]+tmp[1995]*kernel[4]+tmp[1996]*kernel[5]+tmp[2094]*kernel[6]+tmp[2095]*kernel[7]+tmp[2096]*kernel[8];
				ans[1996]<=tmp[1895]*kernel[0]+tmp[1896]*kernel[1]+tmp[1897]*kernel[2]+tmp[1995]*kernel[3]+tmp[1996]*kernel[4]+tmp[1997]*kernel[5]+tmp[2095]*kernel[6]+tmp[2096]*kernel[7]+tmp[2097]*kernel[8];
				ans[1997]<=tmp[1896]*kernel[0]+tmp[1897]*kernel[1]+tmp[1898]*kernel[2]+tmp[1996]*kernel[3]+tmp[1997]*kernel[4]+tmp[1998]*kernel[5]+tmp[2096]*kernel[6]+tmp[2097]*kernel[7]+tmp[2098]*kernel[8];
				ans[1998]<=tmp[1897]*kernel[0]+tmp[1898]*kernel[1]+tmp[1899]*kernel[2]+tmp[1997]*kernel[3]+tmp[1998]*kernel[4]+tmp[1999]*kernel[5]+tmp[2097]*kernel[6]+tmp[2098]*kernel[7]+tmp[2099]*kernel[8];
				ans[1999]<=tmp[1898]*kernel[0]+tmp[1899]*kernel[1]+tmp[1998]*kernel[3]+tmp[1999]*kernel[4]+tmp[2098]*kernel[6]+tmp[2099]*kernel[7];
				ans[2000]<=tmp[1900]*kernel[1]+tmp[1901]*kernel[2]+tmp[2000]*kernel[4]+tmp[2001]*kernel[5]+tmp[2100]*kernel[7]+tmp[2101]*kernel[8];
				ans[2001]<=tmp[1900]*kernel[0]+tmp[1901]*kernel[1]+tmp[1902]*kernel[2]+tmp[2000]*kernel[3]+tmp[2001]*kernel[4]+tmp[2002]*kernel[5]+tmp[2100]*kernel[6]+tmp[2101]*kernel[7]+tmp[2102]*kernel[8];
				ans[2002]<=tmp[1901]*kernel[0]+tmp[1902]*kernel[1]+tmp[1903]*kernel[2]+tmp[2001]*kernel[3]+tmp[2002]*kernel[4]+tmp[2003]*kernel[5]+tmp[2101]*kernel[6]+tmp[2102]*kernel[7]+tmp[2103]*kernel[8];
				ans[2003]<=tmp[1902]*kernel[0]+tmp[1903]*kernel[1]+tmp[1904]*kernel[2]+tmp[2002]*kernel[3]+tmp[2003]*kernel[4]+tmp[2004]*kernel[5]+tmp[2102]*kernel[6]+tmp[2103]*kernel[7]+tmp[2104]*kernel[8];
				ans[2004]<=tmp[1903]*kernel[0]+tmp[1904]*kernel[1]+tmp[1905]*kernel[2]+tmp[2003]*kernel[3]+tmp[2004]*kernel[4]+tmp[2005]*kernel[5]+tmp[2103]*kernel[6]+tmp[2104]*kernel[7]+tmp[2105]*kernel[8];
				ans[2005]<=tmp[1904]*kernel[0]+tmp[1905]*kernel[1]+tmp[1906]*kernel[2]+tmp[2004]*kernel[3]+tmp[2005]*kernel[4]+tmp[2006]*kernel[5]+tmp[2104]*kernel[6]+tmp[2105]*kernel[7]+tmp[2106]*kernel[8];
				ans[2006]<=tmp[1905]*kernel[0]+tmp[1906]*kernel[1]+tmp[1907]*kernel[2]+tmp[2005]*kernel[3]+tmp[2006]*kernel[4]+tmp[2007]*kernel[5]+tmp[2105]*kernel[6]+tmp[2106]*kernel[7]+tmp[2107]*kernel[8];
				ans[2007]<=tmp[1906]*kernel[0]+tmp[1907]*kernel[1]+tmp[1908]*kernel[2]+tmp[2006]*kernel[3]+tmp[2007]*kernel[4]+tmp[2008]*kernel[5]+tmp[2106]*kernel[6]+tmp[2107]*kernel[7]+tmp[2108]*kernel[8];
				ans[2008]<=tmp[1907]*kernel[0]+tmp[1908]*kernel[1]+tmp[1909]*kernel[2]+tmp[2007]*kernel[3]+tmp[2008]*kernel[4]+tmp[2009]*kernel[5]+tmp[2107]*kernel[6]+tmp[2108]*kernel[7]+tmp[2109]*kernel[8];
				ans[2009]<=tmp[1908]*kernel[0]+tmp[1909]*kernel[1]+tmp[1910]*kernel[2]+tmp[2008]*kernel[3]+tmp[2009]*kernel[4]+tmp[2010]*kernel[5]+tmp[2108]*kernel[6]+tmp[2109]*kernel[7]+tmp[2110]*kernel[8];
				ans[2010]<=tmp[1909]*kernel[0]+tmp[1910]*kernel[1]+tmp[1911]*kernel[2]+tmp[2009]*kernel[3]+tmp[2010]*kernel[4]+tmp[2011]*kernel[5]+tmp[2109]*kernel[6]+tmp[2110]*kernel[7]+tmp[2111]*kernel[8];
				ans[2011]<=tmp[1910]*kernel[0]+tmp[1911]*kernel[1]+tmp[1912]*kernel[2]+tmp[2010]*kernel[3]+tmp[2011]*kernel[4]+tmp[2012]*kernel[5]+tmp[2110]*kernel[6]+tmp[2111]*kernel[7]+tmp[2112]*kernel[8];
				ans[2012]<=tmp[1911]*kernel[0]+tmp[1912]*kernel[1]+tmp[1913]*kernel[2]+tmp[2011]*kernel[3]+tmp[2012]*kernel[4]+tmp[2013]*kernel[5]+tmp[2111]*kernel[6]+tmp[2112]*kernel[7]+tmp[2113]*kernel[8];
				ans[2013]<=tmp[1912]*kernel[0]+tmp[1913]*kernel[1]+tmp[1914]*kernel[2]+tmp[2012]*kernel[3]+tmp[2013]*kernel[4]+tmp[2014]*kernel[5]+tmp[2112]*kernel[6]+tmp[2113]*kernel[7]+tmp[2114]*kernel[8];
				ans[2014]<=tmp[1913]*kernel[0]+tmp[1914]*kernel[1]+tmp[1915]*kernel[2]+tmp[2013]*kernel[3]+tmp[2014]*kernel[4]+tmp[2015]*kernel[5]+tmp[2113]*kernel[6]+tmp[2114]*kernel[7]+tmp[2115]*kernel[8];
				ans[2015]<=tmp[1914]*kernel[0]+tmp[1915]*kernel[1]+tmp[1916]*kernel[2]+tmp[2014]*kernel[3]+tmp[2015]*kernel[4]+tmp[2016]*kernel[5]+tmp[2114]*kernel[6]+tmp[2115]*kernel[7]+tmp[2116]*kernel[8];
				ans[2016]<=tmp[1915]*kernel[0]+tmp[1916]*kernel[1]+tmp[1917]*kernel[2]+tmp[2015]*kernel[3]+tmp[2016]*kernel[4]+tmp[2017]*kernel[5]+tmp[2115]*kernel[6]+tmp[2116]*kernel[7]+tmp[2117]*kernel[8];
				ans[2017]<=tmp[1916]*kernel[0]+tmp[1917]*kernel[1]+tmp[1918]*kernel[2]+tmp[2016]*kernel[3]+tmp[2017]*kernel[4]+tmp[2018]*kernel[5]+tmp[2116]*kernel[6]+tmp[2117]*kernel[7]+tmp[2118]*kernel[8];
				ans[2018]<=tmp[1917]*kernel[0]+tmp[1918]*kernel[1]+tmp[1919]*kernel[2]+tmp[2017]*kernel[3]+tmp[2018]*kernel[4]+tmp[2019]*kernel[5]+tmp[2117]*kernel[6]+tmp[2118]*kernel[7]+tmp[2119]*kernel[8];
				ans[2019]<=tmp[1918]*kernel[0]+tmp[1919]*kernel[1]+tmp[1920]*kernel[2]+tmp[2018]*kernel[3]+tmp[2019]*kernel[4]+tmp[2020]*kernel[5]+tmp[2118]*kernel[6]+tmp[2119]*kernel[7]+tmp[2120]*kernel[8];
				ans[2020]<=tmp[1919]*kernel[0]+tmp[1920]*kernel[1]+tmp[1921]*kernel[2]+tmp[2019]*kernel[3]+tmp[2020]*kernel[4]+tmp[2021]*kernel[5]+tmp[2119]*kernel[6]+tmp[2120]*kernel[7]+tmp[2121]*kernel[8];
				ans[2021]<=tmp[1920]*kernel[0]+tmp[1921]*kernel[1]+tmp[1922]*kernel[2]+tmp[2020]*kernel[3]+tmp[2021]*kernel[4]+tmp[2022]*kernel[5]+tmp[2120]*kernel[6]+tmp[2121]*kernel[7]+tmp[2122]*kernel[8];
				ans[2022]<=tmp[1921]*kernel[0]+tmp[1922]*kernel[1]+tmp[1923]*kernel[2]+tmp[2021]*kernel[3]+tmp[2022]*kernel[4]+tmp[2023]*kernel[5]+tmp[2121]*kernel[6]+tmp[2122]*kernel[7]+tmp[2123]*kernel[8];
				ans[2023]<=tmp[1922]*kernel[0]+tmp[1923]*kernel[1]+tmp[1924]*kernel[2]+tmp[2022]*kernel[3]+tmp[2023]*kernel[4]+tmp[2024]*kernel[5]+tmp[2122]*kernel[6]+tmp[2123]*kernel[7]+tmp[2124]*kernel[8];
				ans[2024]<=tmp[1923]*kernel[0]+tmp[1924]*kernel[1]+tmp[1925]*kernel[2]+tmp[2023]*kernel[3]+tmp[2024]*kernel[4]+tmp[2025]*kernel[5]+tmp[2123]*kernel[6]+tmp[2124]*kernel[7]+tmp[2125]*kernel[8];
				ans[2025]<=tmp[1924]*kernel[0]+tmp[1925]*kernel[1]+tmp[1926]*kernel[2]+tmp[2024]*kernel[3]+tmp[2025]*kernel[4]+tmp[2026]*kernel[5]+tmp[2124]*kernel[6]+tmp[2125]*kernel[7]+tmp[2126]*kernel[8];
				ans[2026]<=tmp[1925]*kernel[0]+tmp[1926]*kernel[1]+tmp[1927]*kernel[2]+tmp[2025]*kernel[3]+tmp[2026]*kernel[4]+tmp[2027]*kernel[5]+tmp[2125]*kernel[6]+tmp[2126]*kernel[7]+tmp[2127]*kernel[8];
				ans[2027]<=tmp[1926]*kernel[0]+tmp[1927]*kernel[1]+tmp[1928]*kernel[2]+tmp[2026]*kernel[3]+tmp[2027]*kernel[4]+tmp[2028]*kernel[5]+tmp[2126]*kernel[6]+tmp[2127]*kernel[7]+tmp[2128]*kernel[8];
				ans[2028]<=tmp[1927]*kernel[0]+tmp[1928]*kernel[1]+tmp[1929]*kernel[2]+tmp[2027]*kernel[3]+tmp[2028]*kernel[4]+tmp[2029]*kernel[5]+tmp[2127]*kernel[6]+tmp[2128]*kernel[7]+tmp[2129]*kernel[8];
				ans[2029]<=tmp[1928]*kernel[0]+tmp[1929]*kernel[1]+tmp[1930]*kernel[2]+tmp[2028]*kernel[3]+tmp[2029]*kernel[4]+tmp[2030]*kernel[5]+tmp[2128]*kernel[6]+tmp[2129]*kernel[7]+tmp[2130]*kernel[8];
				ans[2030]<=tmp[1929]*kernel[0]+tmp[1930]*kernel[1]+tmp[1931]*kernel[2]+tmp[2029]*kernel[3]+tmp[2030]*kernel[4]+tmp[2031]*kernel[5]+tmp[2129]*kernel[6]+tmp[2130]*kernel[7]+tmp[2131]*kernel[8];
				ans[2031]<=tmp[1930]*kernel[0]+tmp[1931]*kernel[1]+tmp[1932]*kernel[2]+tmp[2030]*kernel[3]+tmp[2031]*kernel[4]+tmp[2032]*kernel[5]+tmp[2130]*kernel[6]+tmp[2131]*kernel[7]+tmp[2132]*kernel[8];
				ans[2032]<=tmp[1931]*kernel[0]+tmp[1932]*kernel[1]+tmp[1933]*kernel[2]+tmp[2031]*kernel[3]+tmp[2032]*kernel[4]+tmp[2033]*kernel[5]+tmp[2131]*kernel[6]+tmp[2132]*kernel[7]+tmp[2133]*kernel[8];
				ans[2033]<=tmp[1932]*kernel[0]+tmp[1933]*kernel[1]+tmp[1934]*kernel[2]+tmp[2032]*kernel[3]+tmp[2033]*kernel[4]+tmp[2034]*kernel[5]+tmp[2132]*kernel[6]+tmp[2133]*kernel[7]+tmp[2134]*kernel[8];
				ans[2034]<=tmp[1933]*kernel[0]+tmp[1934]*kernel[1]+tmp[1935]*kernel[2]+tmp[2033]*kernel[3]+tmp[2034]*kernel[4]+tmp[2035]*kernel[5]+tmp[2133]*kernel[6]+tmp[2134]*kernel[7]+tmp[2135]*kernel[8];
				ans[2035]<=tmp[1934]*kernel[0]+tmp[1935]*kernel[1]+tmp[1936]*kernel[2]+tmp[2034]*kernel[3]+tmp[2035]*kernel[4]+tmp[2036]*kernel[5]+tmp[2134]*kernel[6]+tmp[2135]*kernel[7]+tmp[2136]*kernel[8];
				ans[2036]<=tmp[1935]*kernel[0]+tmp[1936]*kernel[1]+tmp[1937]*kernel[2]+tmp[2035]*kernel[3]+tmp[2036]*kernel[4]+tmp[2037]*kernel[5]+tmp[2135]*kernel[6]+tmp[2136]*kernel[7]+tmp[2137]*kernel[8];
				ans[2037]<=tmp[1936]*kernel[0]+tmp[1937]*kernel[1]+tmp[1938]*kernel[2]+tmp[2036]*kernel[3]+tmp[2037]*kernel[4]+tmp[2038]*kernel[5]+tmp[2136]*kernel[6]+tmp[2137]*kernel[7]+tmp[2138]*kernel[8];
				ans[2038]<=tmp[1937]*kernel[0]+tmp[1938]*kernel[1]+tmp[1939]*kernel[2]+tmp[2037]*kernel[3]+tmp[2038]*kernel[4]+tmp[2039]*kernel[5]+tmp[2137]*kernel[6]+tmp[2138]*kernel[7]+tmp[2139]*kernel[8];
				ans[2039]<=tmp[1938]*kernel[0]+tmp[1939]*kernel[1]+tmp[1940]*kernel[2]+tmp[2038]*kernel[3]+tmp[2039]*kernel[4]+tmp[2040]*kernel[5]+tmp[2138]*kernel[6]+tmp[2139]*kernel[7]+tmp[2140]*kernel[8];
				ans[2040]<=tmp[1939]*kernel[0]+tmp[1940]*kernel[1]+tmp[1941]*kernel[2]+tmp[2039]*kernel[3]+tmp[2040]*kernel[4]+tmp[2041]*kernel[5]+tmp[2139]*kernel[6]+tmp[2140]*kernel[7]+tmp[2141]*kernel[8];
				ans[2041]<=tmp[1940]*kernel[0]+tmp[1941]*kernel[1]+tmp[1942]*kernel[2]+tmp[2040]*kernel[3]+tmp[2041]*kernel[4]+tmp[2042]*kernel[5]+tmp[2140]*kernel[6]+tmp[2141]*kernel[7]+tmp[2142]*kernel[8];
				ans[2042]<=tmp[1941]*kernel[0]+tmp[1942]*kernel[1]+tmp[1943]*kernel[2]+tmp[2041]*kernel[3]+tmp[2042]*kernel[4]+tmp[2043]*kernel[5]+tmp[2141]*kernel[6]+tmp[2142]*kernel[7]+tmp[2143]*kernel[8];
				ans[2043]<=tmp[1942]*kernel[0]+tmp[1943]*kernel[1]+tmp[1944]*kernel[2]+tmp[2042]*kernel[3]+tmp[2043]*kernel[4]+tmp[2044]*kernel[5]+tmp[2142]*kernel[6]+tmp[2143]*kernel[7]+tmp[2144]*kernel[8];
				ans[2044]<=tmp[1943]*kernel[0]+tmp[1944]*kernel[1]+tmp[1945]*kernel[2]+tmp[2043]*kernel[3]+tmp[2044]*kernel[4]+tmp[2045]*kernel[5]+tmp[2143]*kernel[6]+tmp[2144]*kernel[7]+tmp[2145]*kernel[8];
				ans[2045]<=tmp[1944]*kernel[0]+tmp[1945]*kernel[1]+tmp[1946]*kernel[2]+tmp[2044]*kernel[3]+tmp[2045]*kernel[4]+tmp[2046]*kernel[5]+tmp[2144]*kernel[6]+tmp[2145]*kernel[7]+tmp[2146]*kernel[8];
				ans[2046]<=tmp[1945]*kernel[0]+tmp[1946]*kernel[1]+tmp[1947]*kernel[2]+tmp[2045]*kernel[3]+tmp[2046]*kernel[4]+tmp[2047]*kernel[5]+tmp[2145]*kernel[6]+tmp[2146]*kernel[7]+tmp[2147]*kernel[8];
				ans[2047]<=tmp[1946]*kernel[0]+tmp[1947]*kernel[1]+tmp[1948]*kernel[2]+tmp[2046]*kernel[3]+tmp[2047]*kernel[4]+tmp[2048]*kernel[5]+tmp[2146]*kernel[6]+tmp[2147]*kernel[7]+tmp[2148]*kernel[8];
				ans[2048]<=tmp[1947]*kernel[0]+tmp[1948]*kernel[1]+tmp[1949]*kernel[2]+tmp[2047]*kernel[3]+tmp[2048]*kernel[4]+tmp[2049]*kernel[5]+tmp[2147]*kernel[6]+tmp[2148]*kernel[7]+tmp[2149]*kernel[8];
				ans[2049]<=tmp[1948]*kernel[0]+tmp[1949]*kernel[1]+tmp[1950]*kernel[2]+tmp[2048]*kernel[3]+tmp[2049]*kernel[4]+tmp[2050]*kernel[5]+tmp[2148]*kernel[6]+tmp[2149]*kernel[7]+tmp[2150]*kernel[8];
				ans[2050]<=tmp[1949]*kernel[0]+tmp[1950]*kernel[1]+tmp[1951]*kernel[2]+tmp[2049]*kernel[3]+tmp[2050]*kernel[4]+tmp[2051]*kernel[5]+tmp[2149]*kernel[6]+tmp[2150]*kernel[7]+tmp[2151]*kernel[8];
				ans[2051]<=tmp[1950]*kernel[0]+tmp[1951]*kernel[1]+tmp[1952]*kernel[2]+tmp[2050]*kernel[3]+tmp[2051]*kernel[4]+tmp[2052]*kernel[5]+tmp[2150]*kernel[6]+tmp[2151]*kernel[7]+tmp[2152]*kernel[8];
				ans[2052]<=tmp[1951]*kernel[0]+tmp[1952]*kernel[1]+tmp[1953]*kernel[2]+tmp[2051]*kernel[3]+tmp[2052]*kernel[4]+tmp[2053]*kernel[5]+tmp[2151]*kernel[6]+tmp[2152]*kernel[7]+tmp[2153]*kernel[8];
				ans[2053]<=tmp[1952]*kernel[0]+tmp[1953]*kernel[1]+tmp[1954]*kernel[2]+tmp[2052]*kernel[3]+tmp[2053]*kernel[4]+tmp[2054]*kernel[5]+tmp[2152]*kernel[6]+tmp[2153]*kernel[7]+tmp[2154]*kernel[8];
				ans[2054]<=tmp[1953]*kernel[0]+tmp[1954]*kernel[1]+tmp[1955]*kernel[2]+tmp[2053]*kernel[3]+tmp[2054]*kernel[4]+tmp[2055]*kernel[5]+tmp[2153]*kernel[6]+tmp[2154]*kernel[7]+tmp[2155]*kernel[8];
				ans[2055]<=tmp[1954]*kernel[0]+tmp[1955]*kernel[1]+tmp[1956]*kernel[2]+tmp[2054]*kernel[3]+tmp[2055]*kernel[4]+tmp[2056]*kernel[5]+tmp[2154]*kernel[6]+tmp[2155]*kernel[7]+tmp[2156]*kernel[8];
				ans[2056]<=tmp[1955]*kernel[0]+tmp[1956]*kernel[1]+tmp[1957]*kernel[2]+tmp[2055]*kernel[3]+tmp[2056]*kernel[4]+tmp[2057]*kernel[5]+tmp[2155]*kernel[6]+tmp[2156]*kernel[7]+tmp[2157]*kernel[8];
				ans[2057]<=tmp[1956]*kernel[0]+tmp[1957]*kernel[1]+tmp[1958]*kernel[2]+tmp[2056]*kernel[3]+tmp[2057]*kernel[4]+tmp[2058]*kernel[5]+tmp[2156]*kernel[6]+tmp[2157]*kernel[7]+tmp[2158]*kernel[8];
				ans[2058]<=tmp[1957]*kernel[0]+tmp[1958]*kernel[1]+tmp[1959]*kernel[2]+tmp[2057]*kernel[3]+tmp[2058]*kernel[4]+tmp[2059]*kernel[5]+tmp[2157]*kernel[6]+tmp[2158]*kernel[7]+tmp[2159]*kernel[8];
				ans[2059]<=tmp[1958]*kernel[0]+tmp[1959]*kernel[1]+tmp[1960]*kernel[2]+tmp[2058]*kernel[3]+tmp[2059]*kernel[4]+tmp[2060]*kernel[5]+tmp[2158]*kernel[6]+tmp[2159]*kernel[7]+tmp[2160]*kernel[8];
				ans[2060]<=tmp[1959]*kernel[0]+tmp[1960]*kernel[1]+tmp[1961]*kernel[2]+tmp[2059]*kernel[3]+tmp[2060]*kernel[4]+tmp[2061]*kernel[5]+tmp[2159]*kernel[6]+tmp[2160]*kernel[7]+tmp[2161]*kernel[8];
				ans[2061]<=tmp[1960]*kernel[0]+tmp[1961]*kernel[1]+tmp[1962]*kernel[2]+tmp[2060]*kernel[3]+tmp[2061]*kernel[4]+tmp[2062]*kernel[5]+tmp[2160]*kernel[6]+tmp[2161]*kernel[7]+tmp[2162]*kernel[8];
				ans[2062]<=tmp[1961]*kernel[0]+tmp[1962]*kernel[1]+tmp[1963]*kernel[2]+tmp[2061]*kernel[3]+tmp[2062]*kernel[4]+tmp[2063]*kernel[5]+tmp[2161]*kernel[6]+tmp[2162]*kernel[7]+tmp[2163]*kernel[8];
				ans[2063]<=tmp[1962]*kernel[0]+tmp[1963]*kernel[1]+tmp[1964]*kernel[2]+tmp[2062]*kernel[3]+tmp[2063]*kernel[4]+tmp[2064]*kernel[5]+tmp[2162]*kernel[6]+tmp[2163]*kernel[7]+tmp[2164]*kernel[8];
				ans[2064]<=tmp[1963]*kernel[0]+tmp[1964]*kernel[1]+tmp[1965]*kernel[2]+tmp[2063]*kernel[3]+tmp[2064]*kernel[4]+tmp[2065]*kernel[5]+tmp[2163]*kernel[6]+tmp[2164]*kernel[7]+tmp[2165]*kernel[8];
				ans[2065]<=tmp[1964]*kernel[0]+tmp[1965]*kernel[1]+tmp[1966]*kernel[2]+tmp[2064]*kernel[3]+tmp[2065]*kernel[4]+tmp[2066]*kernel[5]+tmp[2164]*kernel[6]+tmp[2165]*kernel[7]+tmp[2166]*kernel[8];
				ans[2066]<=tmp[1965]*kernel[0]+tmp[1966]*kernel[1]+tmp[1967]*kernel[2]+tmp[2065]*kernel[3]+tmp[2066]*kernel[4]+tmp[2067]*kernel[5]+tmp[2165]*kernel[6]+tmp[2166]*kernel[7]+tmp[2167]*kernel[8];
				ans[2067]<=tmp[1966]*kernel[0]+tmp[1967]*kernel[1]+tmp[1968]*kernel[2]+tmp[2066]*kernel[3]+tmp[2067]*kernel[4]+tmp[2068]*kernel[5]+tmp[2166]*kernel[6]+tmp[2167]*kernel[7]+tmp[2168]*kernel[8];
				ans[2068]<=tmp[1967]*kernel[0]+tmp[1968]*kernel[1]+tmp[1969]*kernel[2]+tmp[2067]*kernel[3]+tmp[2068]*kernel[4]+tmp[2069]*kernel[5]+tmp[2167]*kernel[6]+tmp[2168]*kernel[7]+tmp[2169]*kernel[8];
				ans[2069]<=tmp[1968]*kernel[0]+tmp[1969]*kernel[1]+tmp[1970]*kernel[2]+tmp[2068]*kernel[3]+tmp[2069]*kernel[4]+tmp[2070]*kernel[5]+tmp[2168]*kernel[6]+tmp[2169]*kernel[7]+tmp[2170]*kernel[8];
				ans[2070]<=tmp[1969]*kernel[0]+tmp[1970]*kernel[1]+tmp[1971]*kernel[2]+tmp[2069]*kernel[3]+tmp[2070]*kernel[4]+tmp[2071]*kernel[5]+tmp[2169]*kernel[6]+tmp[2170]*kernel[7]+tmp[2171]*kernel[8];
				ans[2071]<=tmp[1970]*kernel[0]+tmp[1971]*kernel[1]+tmp[1972]*kernel[2]+tmp[2070]*kernel[3]+tmp[2071]*kernel[4]+tmp[2072]*kernel[5]+tmp[2170]*kernel[6]+tmp[2171]*kernel[7]+tmp[2172]*kernel[8];
				ans[2072]<=tmp[1971]*kernel[0]+tmp[1972]*kernel[1]+tmp[1973]*kernel[2]+tmp[2071]*kernel[3]+tmp[2072]*kernel[4]+tmp[2073]*kernel[5]+tmp[2171]*kernel[6]+tmp[2172]*kernel[7]+tmp[2173]*kernel[8];
				ans[2073]<=tmp[1972]*kernel[0]+tmp[1973]*kernel[1]+tmp[1974]*kernel[2]+tmp[2072]*kernel[3]+tmp[2073]*kernel[4]+tmp[2074]*kernel[5]+tmp[2172]*kernel[6]+tmp[2173]*kernel[7]+tmp[2174]*kernel[8];
				ans[2074]<=tmp[1973]*kernel[0]+tmp[1974]*kernel[1]+tmp[1975]*kernel[2]+tmp[2073]*kernel[3]+tmp[2074]*kernel[4]+tmp[2075]*kernel[5]+tmp[2173]*kernel[6]+tmp[2174]*kernel[7]+tmp[2175]*kernel[8];
				ans[2075]<=tmp[1974]*kernel[0]+tmp[1975]*kernel[1]+tmp[1976]*kernel[2]+tmp[2074]*kernel[3]+tmp[2075]*kernel[4]+tmp[2076]*kernel[5]+tmp[2174]*kernel[6]+tmp[2175]*kernel[7]+tmp[2176]*kernel[8];
				ans[2076]<=tmp[1975]*kernel[0]+tmp[1976]*kernel[1]+tmp[1977]*kernel[2]+tmp[2075]*kernel[3]+tmp[2076]*kernel[4]+tmp[2077]*kernel[5]+tmp[2175]*kernel[6]+tmp[2176]*kernel[7]+tmp[2177]*kernel[8];
				ans[2077]<=tmp[1976]*kernel[0]+tmp[1977]*kernel[1]+tmp[1978]*kernel[2]+tmp[2076]*kernel[3]+tmp[2077]*kernel[4]+tmp[2078]*kernel[5]+tmp[2176]*kernel[6]+tmp[2177]*kernel[7]+tmp[2178]*kernel[8];
				ans[2078]<=tmp[1977]*kernel[0]+tmp[1978]*kernel[1]+tmp[1979]*kernel[2]+tmp[2077]*kernel[3]+tmp[2078]*kernel[4]+tmp[2079]*kernel[5]+tmp[2177]*kernel[6]+tmp[2178]*kernel[7]+tmp[2179]*kernel[8];
				ans[2079]<=tmp[1978]*kernel[0]+tmp[1979]*kernel[1]+tmp[1980]*kernel[2]+tmp[2078]*kernel[3]+tmp[2079]*kernel[4]+tmp[2080]*kernel[5]+tmp[2178]*kernel[6]+tmp[2179]*kernel[7]+tmp[2180]*kernel[8];
				ans[2080]<=tmp[1979]*kernel[0]+tmp[1980]*kernel[1]+tmp[1981]*kernel[2]+tmp[2079]*kernel[3]+tmp[2080]*kernel[4]+tmp[2081]*kernel[5]+tmp[2179]*kernel[6]+tmp[2180]*kernel[7]+tmp[2181]*kernel[8];
				ans[2081]<=tmp[1980]*kernel[0]+tmp[1981]*kernel[1]+tmp[1982]*kernel[2]+tmp[2080]*kernel[3]+tmp[2081]*kernel[4]+tmp[2082]*kernel[5]+tmp[2180]*kernel[6]+tmp[2181]*kernel[7]+tmp[2182]*kernel[8];
				ans[2082]<=tmp[1981]*kernel[0]+tmp[1982]*kernel[1]+tmp[1983]*kernel[2]+tmp[2081]*kernel[3]+tmp[2082]*kernel[4]+tmp[2083]*kernel[5]+tmp[2181]*kernel[6]+tmp[2182]*kernel[7]+tmp[2183]*kernel[8];
				ans[2083]<=tmp[1982]*kernel[0]+tmp[1983]*kernel[1]+tmp[1984]*kernel[2]+tmp[2082]*kernel[3]+tmp[2083]*kernel[4]+tmp[2084]*kernel[5]+tmp[2182]*kernel[6]+tmp[2183]*kernel[7]+tmp[2184]*kernel[8];
				ans[2084]<=tmp[1983]*kernel[0]+tmp[1984]*kernel[1]+tmp[1985]*kernel[2]+tmp[2083]*kernel[3]+tmp[2084]*kernel[4]+tmp[2085]*kernel[5]+tmp[2183]*kernel[6]+tmp[2184]*kernel[7]+tmp[2185]*kernel[8];
				ans[2085]<=tmp[1984]*kernel[0]+tmp[1985]*kernel[1]+tmp[1986]*kernel[2]+tmp[2084]*kernel[3]+tmp[2085]*kernel[4]+tmp[2086]*kernel[5]+tmp[2184]*kernel[6]+tmp[2185]*kernel[7]+tmp[2186]*kernel[8];
				ans[2086]<=tmp[1985]*kernel[0]+tmp[1986]*kernel[1]+tmp[1987]*kernel[2]+tmp[2085]*kernel[3]+tmp[2086]*kernel[4]+tmp[2087]*kernel[5]+tmp[2185]*kernel[6]+tmp[2186]*kernel[7]+tmp[2187]*kernel[8];
				ans[2087]<=tmp[1986]*kernel[0]+tmp[1987]*kernel[1]+tmp[1988]*kernel[2]+tmp[2086]*kernel[3]+tmp[2087]*kernel[4]+tmp[2088]*kernel[5]+tmp[2186]*kernel[6]+tmp[2187]*kernel[7]+tmp[2188]*kernel[8];
				ans[2088]<=tmp[1987]*kernel[0]+tmp[1988]*kernel[1]+tmp[1989]*kernel[2]+tmp[2087]*kernel[3]+tmp[2088]*kernel[4]+tmp[2089]*kernel[5]+tmp[2187]*kernel[6]+tmp[2188]*kernel[7]+tmp[2189]*kernel[8];
				ans[2089]<=tmp[1988]*kernel[0]+tmp[1989]*kernel[1]+tmp[1990]*kernel[2]+tmp[2088]*kernel[3]+tmp[2089]*kernel[4]+tmp[2090]*kernel[5]+tmp[2188]*kernel[6]+tmp[2189]*kernel[7]+tmp[2190]*kernel[8];
				ans[2090]<=tmp[1989]*kernel[0]+tmp[1990]*kernel[1]+tmp[1991]*kernel[2]+tmp[2089]*kernel[3]+tmp[2090]*kernel[4]+tmp[2091]*kernel[5]+tmp[2189]*kernel[6]+tmp[2190]*kernel[7]+tmp[2191]*kernel[8];
				ans[2091]<=tmp[1990]*kernel[0]+tmp[1991]*kernel[1]+tmp[1992]*kernel[2]+tmp[2090]*kernel[3]+tmp[2091]*kernel[4]+tmp[2092]*kernel[5]+tmp[2190]*kernel[6]+tmp[2191]*kernel[7]+tmp[2192]*kernel[8];
				ans[2092]<=tmp[1991]*kernel[0]+tmp[1992]*kernel[1]+tmp[1993]*kernel[2]+tmp[2091]*kernel[3]+tmp[2092]*kernel[4]+tmp[2093]*kernel[5]+tmp[2191]*kernel[6]+tmp[2192]*kernel[7]+tmp[2193]*kernel[8];
				ans[2093]<=tmp[1992]*kernel[0]+tmp[1993]*kernel[1]+tmp[1994]*kernel[2]+tmp[2092]*kernel[3]+tmp[2093]*kernel[4]+tmp[2094]*kernel[5]+tmp[2192]*kernel[6]+tmp[2193]*kernel[7]+tmp[2194]*kernel[8];
				ans[2094]<=tmp[1993]*kernel[0]+tmp[1994]*kernel[1]+tmp[1995]*kernel[2]+tmp[2093]*kernel[3]+tmp[2094]*kernel[4]+tmp[2095]*kernel[5]+tmp[2193]*kernel[6]+tmp[2194]*kernel[7]+tmp[2195]*kernel[8];
				ans[2095]<=tmp[1994]*kernel[0]+tmp[1995]*kernel[1]+tmp[1996]*kernel[2]+tmp[2094]*kernel[3]+tmp[2095]*kernel[4]+tmp[2096]*kernel[5]+tmp[2194]*kernel[6]+tmp[2195]*kernel[7]+tmp[2196]*kernel[8];
				ans[2096]<=tmp[1995]*kernel[0]+tmp[1996]*kernel[1]+tmp[1997]*kernel[2]+tmp[2095]*kernel[3]+tmp[2096]*kernel[4]+tmp[2097]*kernel[5]+tmp[2195]*kernel[6]+tmp[2196]*kernel[7]+tmp[2197]*kernel[8];
				ans[2097]<=tmp[1996]*kernel[0]+tmp[1997]*kernel[1]+tmp[1998]*kernel[2]+tmp[2096]*kernel[3]+tmp[2097]*kernel[4]+tmp[2098]*kernel[5]+tmp[2196]*kernel[6]+tmp[2197]*kernel[7]+tmp[2198]*kernel[8];
				ans[2098]<=tmp[1997]*kernel[0]+tmp[1998]*kernel[1]+tmp[1999]*kernel[2]+tmp[2097]*kernel[3]+tmp[2098]*kernel[4]+tmp[2099]*kernel[5]+tmp[2197]*kernel[6]+tmp[2198]*kernel[7]+tmp[2199]*kernel[8];
				ans[2099]<=tmp[1998]*kernel[0]+tmp[1999]*kernel[1]+tmp[2098]*kernel[3]+tmp[2099]*kernel[4]+tmp[2198]*kernel[6]+tmp[2199]*kernel[7];
				ans[2100]<=tmp[2000]*kernel[1]+tmp[2001]*kernel[2]+tmp[2100]*kernel[4]+tmp[2101]*kernel[5]+tmp[2200]*kernel[7]+tmp[2201]*kernel[8];
				ans[2101]<=tmp[2000]*kernel[0]+tmp[2001]*kernel[1]+tmp[2002]*kernel[2]+tmp[2100]*kernel[3]+tmp[2101]*kernel[4]+tmp[2102]*kernel[5]+tmp[2200]*kernel[6]+tmp[2201]*kernel[7]+tmp[2202]*kernel[8];
				ans[2102]<=tmp[2001]*kernel[0]+tmp[2002]*kernel[1]+tmp[2003]*kernel[2]+tmp[2101]*kernel[3]+tmp[2102]*kernel[4]+tmp[2103]*kernel[5]+tmp[2201]*kernel[6]+tmp[2202]*kernel[7]+tmp[2203]*kernel[8];
				ans[2103]<=tmp[2002]*kernel[0]+tmp[2003]*kernel[1]+tmp[2004]*kernel[2]+tmp[2102]*kernel[3]+tmp[2103]*kernel[4]+tmp[2104]*kernel[5]+tmp[2202]*kernel[6]+tmp[2203]*kernel[7]+tmp[2204]*kernel[8];
				ans[2104]<=tmp[2003]*kernel[0]+tmp[2004]*kernel[1]+tmp[2005]*kernel[2]+tmp[2103]*kernel[3]+tmp[2104]*kernel[4]+tmp[2105]*kernel[5]+tmp[2203]*kernel[6]+tmp[2204]*kernel[7]+tmp[2205]*kernel[8];
				ans[2105]<=tmp[2004]*kernel[0]+tmp[2005]*kernel[1]+tmp[2006]*kernel[2]+tmp[2104]*kernel[3]+tmp[2105]*kernel[4]+tmp[2106]*kernel[5]+tmp[2204]*kernel[6]+tmp[2205]*kernel[7]+tmp[2206]*kernel[8];
				ans[2106]<=tmp[2005]*kernel[0]+tmp[2006]*kernel[1]+tmp[2007]*kernel[2]+tmp[2105]*kernel[3]+tmp[2106]*kernel[4]+tmp[2107]*kernel[5]+tmp[2205]*kernel[6]+tmp[2206]*kernel[7]+tmp[2207]*kernel[8];
				ans[2107]<=tmp[2006]*kernel[0]+tmp[2007]*kernel[1]+tmp[2008]*kernel[2]+tmp[2106]*kernel[3]+tmp[2107]*kernel[4]+tmp[2108]*kernel[5]+tmp[2206]*kernel[6]+tmp[2207]*kernel[7]+tmp[2208]*kernel[8];
				ans[2108]<=tmp[2007]*kernel[0]+tmp[2008]*kernel[1]+tmp[2009]*kernel[2]+tmp[2107]*kernel[3]+tmp[2108]*kernel[4]+tmp[2109]*kernel[5]+tmp[2207]*kernel[6]+tmp[2208]*kernel[7]+tmp[2209]*kernel[8];
				ans[2109]<=tmp[2008]*kernel[0]+tmp[2009]*kernel[1]+tmp[2010]*kernel[2]+tmp[2108]*kernel[3]+tmp[2109]*kernel[4]+tmp[2110]*kernel[5]+tmp[2208]*kernel[6]+tmp[2209]*kernel[7]+tmp[2210]*kernel[8];
				ans[2110]<=tmp[2009]*kernel[0]+tmp[2010]*kernel[1]+tmp[2011]*kernel[2]+tmp[2109]*kernel[3]+tmp[2110]*kernel[4]+tmp[2111]*kernel[5]+tmp[2209]*kernel[6]+tmp[2210]*kernel[7]+tmp[2211]*kernel[8];
				ans[2111]<=tmp[2010]*kernel[0]+tmp[2011]*kernel[1]+tmp[2012]*kernel[2]+tmp[2110]*kernel[3]+tmp[2111]*kernel[4]+tmp[2112]*kernel[5]+tmp[2210]*kernel[6]+tmp[2211]*kernel[7]+tmp[2212]*kernel[8];
				ans[2112]<=tmp[2011]*kernel[0]+tmp[2012]*kernel[1]+tmp[2013]*kernel[2]+tmp[2111]*kernel[3]+tmp[2112]*kernel[4]+tmp[2113]*kernel[5]+tmp[2211]*kernel[6]+tmp[2212]*kernel[7]+tmp[2213]*kernel[8];
				ans[2113]<=tmp[2012]*kernel[0]+tmp[2013]*kernel[1]+tmp[2014]*kernel[2]+tmp[2112]*kernel[3]+tmp[2113]*kernel[4]+tmp[2114]*kernel[5]+tmp[2212]*kernel[6]+tmp[2213]*kernel[7]+tmp[2214]*kernel[8];
				ans[2114]<=tmp[2013]*kernel[0]+tmp[2014]*kernel[1]+tmp[2015]*kernel[2]+tmp[2113]*kernel[3]+tmp[2114]*kernel[4]+tmp[2115]*kernel[5]+tmp[2213]*kernel[6]+tmp[2214]*kernel[7]+tmp[2215]*kernel[8];
				ans[2115]<=tmp[2014]*kernel[0]+tmp[2015]*kernel[1]+tmp[2016]*kernel[2]+tmp[2114]*kernel[3]+tmp[2115]*kernel[4]+tmp[2116]*kernel[5]+tmp[2214]*kernel[6]+tmp[2215]*kernel[7]+tmp[2216]*kernel[8];
				ans[2116]<=tmp[2015]*kernel[0]+tmp[2016]*kernel[1]+tmp[2017]*kernel[2]+tmp[2115]*kernel[3]+tmp[2116]*kernel[4]+tmp[2117]*kernel[5]+tmp[2215]*kernel[6]+tmp[2216]*kernel[7]+tmp[2217]*kernel[8];
				ans[2117]<=tmp[2016]*kernel[0]+tmp[2017]*kernel[1]+tmp[2018]*kernel[2]+tmp[2116]*kernel[3]+tmp[2117]*kernel[4]+tmp[2118]*kernel[5]+tmp[2216]*kernel[6]+tmp[2217]*kernel[7]+tmp[2218]*kernel[8];
				ans[2118]<=tmp[2017]*kernel[0]+tmp[2018]*kernel[1]+tmp[2019]*kernel[2]+tmp[2117]*kernel[3]+tmp[2118]*kernel[4]+tmp[2119]*kernel[5]+tmp[2217]*kernel[6]+tmp[2218]*kernel[7]+tmp[2219]*kernel[8];
				ans[2119]<=tmp[2018]*kernel[0]+tmp[2019]*kernel[1]+tmp[2020]*kernel[2]+tmp[2118]*kernel[3]+tmp[2119]*kernel[4]+tmp[2120]*kernel[5]+tmp[2218]*kernel[6]+tmp[2219]*kernel[7]+tmp[2220]*kernel[8];
				ans[2120]<=tmp[2019]*kernel[0]+tmp[2020]*kernel[1]+tmp[2021]*kernel[2]+tmp[2119]*kernel[3]+tmp[2120]*kernel[4]+tmp[2121]*kernel[5]+tmp[2219]*kernel[6]+tmp[2220]*kernel[7]+tmp[2221]*kernel[8];
				ans[2121]<=tmp[2020]*kernel[0]+tmp[2021]*kernel[1]+tmp[2022]*kernel[2]+tmp[2120]*kernel[3]+tmp[2121]*kernel[4]+tmp[2122]*kernel[5]+tmp[2220]*kernel[6]+tmp[2221]*kernel[7]+tmp[2222]*kernel[8];
				ans[2122]<=tmp[2021]*kernel[0]+tmp[2022]*kernel[1]+tmp[2023]*kernel[2]+tmp[2121]*kernel[3]+tmp[2122]*kernel[4]+tmp[2123]*kernel[5]+tmp[2221]*kernel[6]+tmp[2222]*kernel[7]+tmp[2223]*kernel[8];
				ans[2123]<=tmp[2022]*kernel[0]+tmp[2023]*kernel[1]+tmp[2024]*kernel[2]+tmp[2122]*kernel[3]+tmp[2123]*kernel[4]+tmp[2124]*kernel[5]+tmp[2222]*kernel[6]+tmp[2223]*kernel[7]+tmp[2224]*kernel[8];
				ans[2124]<=tmp[2023]*kernel[0]+tmp[2024]*kernel[1]+tmp[2025]*kernel[2]+tmp[2123]*kernel[3]+tmp[2124]*kernel[4]+tmp[2125]*kernel[5]+tmp[2223]*kernel[6]+tmp[2224]*kernel[7]+tmp[2225]*kernel[8];
				ans[2125]<=tmp[2024]*kernel[0]+tmp[2025]*kernel[1]+tmp[2026]*kernel[2]+tmp[2124]*kernel[3]+tmp[2125]*kernel[4]+tmp[2126]*kernel[5]+tmp[2224]*kernel[6]+tmp[2225]*kernel[7]+tmp[2226]*kernel[8];
				ans[2126]<=tmp[2025]*kernel[0]+tmp[2026]*kernel[1]+tmp[2027]*kernel[2]+tmp[2125]*kernel[3]+tmp[2126]*kernel[4]+tmp[2127]*kernel[5]+tmp[2225]*kernel[6]+tmp[2226]*kernel[7]+tmp[2227]*kernel[8];
				ans[2127]<=tmp[2026]*kernel[0]+tmp[2027]*kernel[1]+tmp[2028]*kernel[2]+tmp[2126]*kernel[3]+tmp[2127]*kernel[4]+tmp[2128]*kernel[5]+tmp[2226]*kernel[6]+tmp[2227]*kernel[7]+tmp[2228]*kernel[8];
				ans[2128]<=tmp[2027]*kernel[0]+tmp[2028]*kernel[1]+tmp[2029]*kernel[2]+tmp[2127]*kernel[3]+tmp[2128]*kernel[4]+tmp[2129]*kernel[5]+tmp[2227]*kernel[6]+tmp[2228]*kernel[7]+tmp[2229]*kernel[8];
				ans[2129]<=tmp[2028]*kernel[0]+tmp[2029]*kernel[1]+tmp[2030]*kernel[2]+tmp[2128]*kernel[3]+tmp[2129]*kernel[4]+tmp[2130]*kernel[5]+tmp[2228]*kernel[6]+tmp[2229]*kernel[7]+tmp[2230]*kernel[8];
				ans[2130]<=tmp[2029]*kernel[0]+tmp[2030]*kernel[1]+tmp[2031]*kernel[2]+tmp[2129]*kernel[3]+tmp[2130]*kernel[4]+tmp[2131]*kernel[5]+tmp[2229]*kernel[6]+tmp[2230]*kernel[7]+tmp[2231]*kernel[8];
				ans[2131]<=tmp[2030]*kernel[0]+tmp[2031]*kernel[1]+tmp[2032]*kernel[2]+tmp[2130]*kernel[3]+tmp[2131]*kernel[4]+tmp[2132]*kernel[5]+tmp[2230]*kernel[6]+tmp[2231]*kernel[7]+tmp[2232]*kernel[8];
				ans[2132]<=tmp[2031]*kernel[0]+tmp[2032]*kernel[1]+tmp[2033]*kernel[2]+tmp[2131]*kernel[3]+tmp[2132]*kernel[4]+tmp[2133]*kernel[5]+tmp[2231]*kernel[6]+tmp[2232]*kernel[7]+tmp[2233]*kernel[8];
				ans[2133]<=tmp[2032]*kernel[0]+tmp[2033]*kernel[1]+tmp[2034]*kernel[2]+tmp[2132]*kernel[3]+tmp[2133]*kernel[4]+tmp[2134]*kernel[5]+tmp[2232]*kernel[6]+tmp[2233]*kernel[7]+tmp[2234]*kernel[8];
				ans[2134]<=tmp[2033]*kernel[0]+tmp[2034]*kernel[1]+tmp[2035]*kernel[2]+tmp[2133]*kernel[3]+tmp[2134]*kernel[4]+tmp[2135]*kernel[5]+tmp[2233]*kernel[6]+tmp[2234]*kernel[7]+tmp[2235]*kernel[8];
				ans[2135]<=tmp[2034]*kernel[0]+tmp[2035]*kernel[1]+tmp[2036]*kernel[2]+tmp[2134]*kernel[3]+tmp[2135]*kernel[4]+tmp[2136]*kernel[5]+tmp[2234]*kernel[6]+tmp[2235]*kernel[7]+tmp[2236]*kernel[8];
				ans[2136]<=tmp[2035]*kernel[0]+tmp[2036]*kernel[1]+tmp[2037]*kernel[2]+tmp[2135]*kernel[3]+tmp[2136]*kernel[4]+tmp[2137]*kernel[5]+tmp[2235]*kernel[6]+tmp[2236]*kernel[7]+tmp[2237]*kernel[8];
				ans[2137]<=tmp[2036]*kernel[0]+tmp[2037]*kernel[1]+tmp[2038]*kernel[2]+tmp[2136]*kernel[3]+tmp[2137]*kernel[4]+tmp[2138]*kernel[5]+tmp[2236]*kernel[6]+tmp[2237]*kernel[7]+tmp[2238]*kernel[8];
				ans[2138]<=tmp[2037]*kernel[0]+tmp[2038]*kernel[1]+tmp[2039]*kernel[2]+tmp[2137]*kernel[3]+tmp[2138]*kernel[4]+tmp[2139]*kernel[5]+tmp[2237]*kernel[6]+tmp[2238]*kernel[7]+tmp[2239]*kernel[8];
				ans[2139]<=tmp[2038]*kernel[0]+tmp[2039]*kernel[1]+tmp[2040]*kernel[2]+tmp[2138]*kernel[3]+tmp[2139]*kernel[4]+tmp[2140]*kernel[5]+tmp[2238]*kernel[6]+tmp[2239]*kernel[7]+tmp[2240]*kernel[8];
				ans[2140]<=tmp[2039]*kernel[0]+tmp[2040]*kernel[1]+tmp[2041]*kernel[2]+tmp[2139]*kernel[3]+tmp[2140]*kernel[4]+tmp[2141]*kernel[5]+tmp[2239]*kernel[6]+tmp[2240]*kernel[7]+tmp[2241]*kernel[8];
				ans[2141]<=tmp[2040]*kernel[0]+tmp[2041]*kernel[1]+tmp[2042]*kernel[2]+tmp[2140]*kernel[3]+tmp[2141]*kernel[4]+tmp[2142]*kernel[5]+tmp[2240]*kernel[6]+tmp[2241]*kernel[7]+tmp[2242]*kernel[8];
				ans[2142]<=tmp[2041]*kernel[0]+tmp[2042]*kernel[1]+tmp[2043]*kernel[2]+tmp[2141]*kernel[3]+tmp[2142]*kernel[4]+tmp[2143]*kernel[5]+tmp[2241]*kernel[6]+tmp[2242]*kernel[7]+tmp[2243]*kernel[8];
				ans[2143]<=tmp[2042]*kernel[0]+tmp[2043]*kernel[1]+tmp[2044]*kernel[2]+tmp[2142]*kernel[3]+tmp[2143]*kernel[4]+tmp[2144]*kernel[5]+tmp[2242]*kernel[6]+tmp[2243]*kernel[7]+tmp[2244]*kernel[8];
				ans[2144]<=tmp[2043]*kernel[0]+tmp[2044]*kernel[1]+tmp[2045]*kernel[2]+tmp[2143]*kernel[3]+tmp[2144]*kernel[4]+tmp[2145]*kernel[5]+tmp[2243]*kernel[6]+tmp[2244]*kernel[7]+tmp[2245]*kernel[8];
				ans[2145]<=tmp[2044]*kernel[0]+tmp[2045]*kernel[1]+tmp[2046]*kernel[2]+tmp[2144]*kernel[3]+tmp[2145]*kernel[4]+tmp[2146]*kernel[5]+tmp[2244]*kernel[6]+tmp[2245]*kernel[7]+tmp[2246]*kernel[8];
				ans[2146]<=tmp[2045]*kernel[0]+tmp[2046]*kernel[1]+tmp[2047]*kernel[2]+tmp[2145]*kernel[3]+tmp[2146]*kernel[4]+tmp[2147]*kernel[5]+tmp[2245]*kernel[6]+tmp[2246]*kernel[7]+tmp[2247]*kernel[8];
				ans[2147]<=tmp[2046]*kernel[0]+tmp[2047]*kernel[1]+tmp[2048]*kernel[2]+tmp[2146]*kernel[3]+tmp[2147]*kernel[4]+tmp[2148]*kernel[5]+tmp[2246]*kernel[6]+tmp[2247]*kernel[7]+tmp[2248]*kernel[8];
				ans[2148]<=tmp[2047]*kernel[0]+tmp[2048]*kernel[1]+tmp[2049]*kernel[2]+tmp[2147]*kernel[3]+tmp[2148]*kernel[4]+tmp[2149]*kernel[5]+tmp[2247]*kernel[6]+tmp[2248]*kernel[7]+tmp[2249]*kernel[8];
				ans[2149]<=tmp[2048]*kernel[0]+tmp[2049]*kernel[1]+tmp[2050]*kernel[2]+tmp[2148]*kernel[3]+tmp[2149]*kernel[4]+tmp[2150]*kernel[5]+tmp[2248]*kernel[6]+tmp[2249]*kernel[7]+tmp[2250]*kernel[8];
				ans[2150]<=tmp[2049]*kernel[0]+tmp[2050]*kernel[1]+tmp[2051]*kernel[2]+tmp[2149]*kernel[3]+tmp[2150]*kernel[4]+tmp[2151]*kernel[5]+tmp[2249]*kernel[6]+tmp[2250]*kernel[7]+tmp[2251]*kernel[8];
				ans[2151]<=tmp[2050]*kernel[0]+tmp[2051]*kernel[1]+tmp[2052]*kernel[2]+tmp[2150]*kernel[3]+tmp[2151]*kernel[4]+tmp[2152]*kernel[5]+tmp[2250]*kernel[6]+tmp[2251]*kernel[7]+tmp[2252]*kernel[8];
				ans[2152]<=tmp[2051]*kernel[0]+tmp[2052]*kernel[1]+tmp[2053]*kernel[2]+tmp[2151]*kernel[3]+tmp[2152]*kernel[4]+tmp[2153]*kernel[5]+tmp[2251]*kernel[6]+tmp[2252]*kernel[7]+tmp[2253]*kernel[8];
				ans[2153]<=tmp[2052]*kernel[0]+tmp[2053]*kernel[1]+tmp[2054]*kernel[2]+tmp[2152]*kernel[3]+tmp[2153]*kernel[4]+tmp[2154]*kernel[5]+tmp[2252]*kernel[6]+tmp[2253]*kernel[7]+tmp[2254]*kernel[8];
				ans[2154]<=tmp[2053]*kernel[0]+tmp[2054]*kernel[1]+tmp[2055]*kernel[2]+tmp[2153]*kernel[3]+tmp[2154]*kernel[4]+tmp[2155]*kernel[5]+tmp[2253]*kernel[6]+tmp[2254]*kernel[7]+tmp[2255]*kernel[8];
				ans[2155]<=tmp[2054]*kernel[0]+tmp[2055]*kernel[1]+tmp[2056]*kernel[2]+tmp[2154]*kernel[3]+tmp[2155]*kernel[4]+tmp[2156]*kernel[5]+tmp[2254]*kernel[6]+tmp[2255]*kernel[7]+tmp[2256]*kernel[8];
				ans[2156]<=tmp[2055]*kernel[0]+tmp[2056]*kernel[1]+tmp[2057]*kernel[2]+tmp[2155]*kernel[3]+tmp[2156]*kernel[4]+tmp[2157]*kernel[5]+tmp[2255]*kernel[6]+tmp[2256]*kernel[7]+tmp[2257]*kernel[8];
				ans[2157]<=tmp[2056]*kernel[0]+tmp[2057]*kernel[1]+tmp[2058]*kernel[2]+tmp[2156]*kernel[3]+tmp[2157]*kernel[4]+tmp[2158]*kernel[5]+tmp[2256]*kernel[6]+tmp[2257]*kernel[7]+tmp[2258]*kernel[8];
				ans[2158]<=tmp[2057]*kernel[0]+tmp[2058]*kernel[1]+tmp[2059]*kernel[2]+tmp[2157]*kernel[3]+tmp[2158]*kernel[4]+tmp[2159]*kernel[5]+tmp[2257]*kernel[6]+tmp[2258]*kernel[7]+tmp[2259]*kernel[8];
				ans[2159]<=tmp[2058]*kernel[0]+tmp[2059]*kernel[1]+tmp[2060]*kernel[2]+tmp[2158]*kernel[3]+tmp[2159]*kernel[4]+tmp[2160]*kernel[5]+tmp[2258]*kernel[6]+tmp[2259]*kernel[7]+tmp[2260]*kernel[8];
				ans[2160]<=tmp[2059]*kernel[0]+tmp[2060]*kernel[1]+tmp[2061]*kernel[2]+tmp[2159]*kernel[3]+tmp[2160]*kernel[4]+tmp[2161]*kernel[5]+tmp[2259]*kernel[6]+tmp[2260]*kernel[7]+tmp[2261]*kernel[8];
				ans[2161]<=tmp[2060]*kernel[0]+tmp[2061]*kernel[1]+tmp[2062]*kernel[2]+tmp[2160]*kernel[3]+tmp[2161]*kernel[4]+tmp[2162]*kernel[5]+tmp[2260]*kernel[6]+tmp[2261]*kernel[7]+tmp[2262]*kernel[8];
				ans[2162]<=tmp[2061]*kernel[0]+tmp[2062]*kernel[1]+tmp[2063]*kernel[2]+tmp[2161]*kernel[3]+tmp[2162]*kernel[4]+tmp[2163]*kernel[5]+tmp[2261]*kernel[6]+tmp[2262]*kernel[7]+tmp[2263]*kernel[8];
				ans[2163]<=tmp[2062]*kernel[0]+tmp[2063]*kernel[1]+tmp[2064]*kernel[2]+tmp[2162]*kernel[3]+tmp[2163]*kernel[4]+tmp[2164]*kernel[5]+tmp[2262]*kernel[6]+tmp[2263]*kernel[7]+tmp[2264]*kernel[8];
				ans[2164]<=tmp[2063]*kernel[0]+tmp[2064]*kernel[1]+tmp[2065]*kernel[2]+tmp[2163]*kernel[3]+tmp[2164]*kernel[4]+tmp[2165]*kernel[5]+tmp[2263]*kernel[6]+tmp[2264]*kernel[7]+tmp[2265]*kernel[8];
				ans[2165]<=tmp[2064]*kernel[0]+tmp[2065]*kernel[1]+tmp[2066]*kernel[2]+tmp[2164]*kernel[3]+tmp[2165]*kernel[4]+tmp[2166]*kernel[5]+tmp[2264]*kernel[6]+tmp[2265]*kernel[7]+tmp[2266]*kernel[8];
				ans[2166]<=tmp[2065]*kernel[0]+tmp[2066]*kernel[1]+tmp[2067]*kernel[2]+tmp[2165]*kernel[3]+tmp[2166]*kernel[4]+tmp[2167]*kernel[5]+tmp[2265]*kernel[6]+tmp[2266]*kernel[7]+tmp[2267]*kernel[8];
				ans[2167]<=tmp[2066]*kernel[0]+tmp[2067]*kernel[1]+tmp[2068]*kernel[2]+tmp[2166]*kernel[3]+tmp[2167]*kernel[4]+tmp[2168]*kernel[5]+tmp[2266]*kernel[6]+tmp[2267]*kernel[7]+tmp[2268]*kernel[8];
				ans[2168]<=tmp[2067]*kernel[0]+tmp[2068]*kernel[1]+tmp[2069]*kernel[2]+tmp[2167]*kernel[3]+tmp[2168]*kernel[4]+tmp[2169]*kernel[5]+tmp[2267]*kernel[6]+tmp[2268]*kernel[7]+tmp[2269]*kernel[8];
				ans[2169]<=tmp[2068]*kernel[0]+tmp[2069]*kernel[1]+tmp[2070]*kernel[2]+tmp[2168]*kernel[3]+tmp[2169]*kernel[4]+tmp[2170]*kernel[5]+tmp[2268]*kernel[6]+tmp[2269]*kernel[7]+tmp[2270]*kernel[8];
				ans[2170]<=tmp[2069]*kernel[0]+tmp[2070]*kernel[1]+tmp[2071]*kernel[2]+tmp[2169]*kernel[3]+tmp[2170]*kernel[4]+tmp[2171]*kernel[5]+tmp[2269]*kernel[6]+tmp[2270]*kernel[7]+tmp[2271]*kernel[8];
				ans[2171]<=tmp[2070]*kernel[0]+tmp[2071]*kernel[1]+tmp[2072]*kernel[2]+tmp[2170]*kernel[3]+tmp[2171]*kernel[4]+tmp[2172]*kernel[5]+tmp[2270]*kernel[6]+tmp[2271]*kernel[7]+tmp[2272]*kernel[8];
				ans[2172]<=tmp[2071]*kernel[0]+tmp[2072]*kernel[1]+tmp[2073]*kernel[2]+tmp[2171]*kernel[3]+tmp[2172]*kernel[4]+tmp[2173]*kernel[5]+tmp[2271]*kernel[6]+tmp[2272]*kernel[7]+tmp[2273]*kernel[8];
				ans[2173]<=tmp[2072]*kernel[0]+tmp[2073]*kernel[1]+tmp[2074]*kernel[2]+tmp[2172]*kernel[3]+tmp[2173]*kernel[4]+tmp[2174]*kernel[5]+tmp[2272]*kernel[6]+tmp[2273]*kernel[7]+tmp[2274]*kernel[8];
				ans[2174]<=tmp[2073]*kernel[0]+tmp[2074]*kernel[1]+tmp[2075]*kernel[2]+tmp[2173]*kernel[3]+tmp[2174]*kernel[4]+tmp[2175]*kernel[5]+tmp[2273]*kernel[6]+tmp[2274]*kernel[7]+tmp[2275]*kernel[8];
				ans[2175]<=tmp[2074]*kernel[0]+tmp[2075]*kernel[1]+tmp[2076]*kernel[2]+tmp[2174]*kernel[3]+tmp[2175]*kernel[4]+tmp[2176]*kernel[5]+tmp[2274]*kernel[6]+tmp[2275]*kernel[7]+tmp[2276]*kernel[8];
				ans[2176]<=tmp[2075]*kernel[0]+tmp[2076]*kernel[1]+tmp[2077]*kernel[2]+tmp[2175]*kernel[3]+tmp[2176]*kernel[4]+tmp[2177]*kernel[5]+tmp[2275]*kernel[6]+tmp[2276]*kernel[7]+tmp[2277]*kernel[8];
				ans[2177]<=tmp[2076]*kernel[0]+tmp[2077]*kernel[1]+tmp[2078]*kernel[2]+tmp[2176]*kernel[3]+tmp[2177]*kernel[4]+tmp[2178]*kernel[5]+tmp[2276]*kernel[6]+tmp[2277]*kernel[7]+tmp[2278]*kernel[8];
				ans[2178]<=tmp[2077]*kernel[0]+tmp[2078]*kernel[1]+tmp[2079]*kernel[2]+tmp[2177]*kernel[3]+tmp[2178]*kernel[4]+tmp[2179]*kernel[5]+tmp[2277]*kernel[6]+tmp[2278]*kernel[7]+tmp[2279]*kernel[8];
				ans[2179]<=tmp[2078]*kernel[0]+tmp[2079]*kernel[1]+tmp[2080]*kernel[2]+tmp[2178]*kernel[3]+tmp[2179]*kernel[4]+tmp[2180]*kernel[5]+tmp[2278]*kernel[6]+tmp[2279]*kernel[7]+tmp[2280]*kernel[8];
				ans[2180]<=tmp[2079]*kernel[0]+tmp[2080]*kernel[1]+tmp[2081]*kernel[2]+tmp[2179]*kernel[3]+tmp[2180]*kernel[4]+tmp[2181]*kernel[5]+tmp[2279]*kernel[6]+tmp[2280]*kernel[7]+tmp[2281]*kernel[8];
				ans[2181]<=tmp[2080]*kernel[0]+tmp[2081]*kernel[1]+tmp[2082]*kernel[2]+tmp[2180]*kernel[3]+tmp[2181]*kernel[4]+tmp[2182]*kernel[5]+tmp[2280]*kernel[6]+tmp[2281]*kernel[7]+tmp[2282]*kernel[8];
				ans[2182]<=tmp[2081]*kernel[0]+tmp[2082]*kernel[1]+tmp[2083]*kernel[2]+tmp[2181]*kernel[3]+tmp[2182]*kernel[4]+tmp[2183]*kernel[5]+tmp[2281]*kernel[6]+tmp[2282]*kernel[7]+tmp[2283]*kernel[8];
				ans[2183]<=tmp[2082]*kernel[0]+tmp[2083]*kernel[1]+tmp[2084]*kernel[2]+tmp[2182]*kernel[3]+tmp[2183]*kernel[4]+tmp[2184]*kernel[5]+tmp[2282]*kernel[6]+tmp[2283]*kernel[7]+tmp[2284]*kernel[8];
				ans[2184]<=tmp[2083]*kernel[0]+tmp[2084]*kernel[1]+tmp[2085]*kernel[2]+tmp[2183]*kernel[3]+tmp[2184]*kernel[4]+tmp[2185]*kernel[5]+tmp[2283]*kernel[6]+tmp[2284]*kernel[7]+tmp[2285]*kernel[8];
				ans[2185]<=tmp[2084]*kernel[0]+tmp[2085]*kernel[1]+tmp[2086]*kernel[2]+tmp[2184]*kernel[3]+tmp[2185]*kernel[4]+tmp[2186]*kernel[5]+tmp[2284]*kernel[6]+tmp[2285]*kernel[7]+tmp[2286]*kernel[8];
				ans[2186]<=tmp[2085]*kernel[0]+tmp[2086]*kernel[1]+tmp[2087]*kernel[2]+tmp[2185]*kernel[3]+tmp[2186]*kernel[4]+tmp[2187]*kernel[5]+tmp[2285]*kernel[6]+tmp[2286]*kernel[7]+tmp[2287]*kernel[8];
				ans[2187]<=tmp[2086]*kernel[0]+tmp[2087]*kernel[1]+tmp[2088]*kernel[2]+tmp[2186]*kernel[3]+tmp[2187]*kernel[4]+tmp[2188]*kernel[5]+tmp[2286]*kernel[6]+tmp[2287]*kernel[7]+tmp[2288]*kernel[8];
				ans[2188]<=tmp[2087]*kernel[0]+tmp[2088]*kernel[1]+tmp[2089]*kernel[2]+tmp[2187]*kernel[3]+tmp[2188]*kernel[4]+tmp[2189]*kernel[5]+tmp[2287]*kernel[6]+tmp[2288]*kernel[7]+tmp[2289]*kernel[8];
				ans[2189]<=tmp[2088]*kernel[0]+tmp[2089]*kernel[1]+tmp[2090]*kernel[2]+tmp[2188]*kernel[3]+tmp[2189]*kernel[4]+tmp[2190]*kernel[5]+tmp[2288]*kernel[6]+tmp[2289]*kernel[7]+tmp[2290]*kernel[8];
				ans[2190]<=tmp[2089]*kernel[0]+tmp[2090]*kernel[1]+tmp[2091]*kernel[2]+tmp[2189]*kernel[3]+tmp[2190]*kernel[4]+tmp[2191]*kernel[5]+tmp[2289]*kernel[6]+tmp[2290]*kernel[7]+tmp[2291]*kernel[8];
				ans[2191]<=tmp[2090]*kernel[0]+tmp[2091]*kernel[1]+tmp[2092]*kernel[2]+tmp[2190]*kernel[3]+tmp[2191]*kernel[4]+tmp[2192]*kernel[5]+tmp[2290]*kernel[6]+tmp[2291]*kernel[7]+tmp[2292]*kernel[8];
				ans[2192]<=tmp[2091]*kernel[0]+tmp[2092]*kernel[1]+tmp[2093]*kernel[2]+tmp[2191]*kernel[3]+tmp[2192]*kernel[4]+tmp[2193]*kernel[5]+tmp[2291]*kernel[6]+tmp[2292]*kernel[7]+tmp[2293]*kernel[8];
				ans[2193]<=tmp[2092]*kernel[0]+tmp[2093]*kernel[1]+tmp[2094]*kernel[2]+tmp[2192]*kernel[3]+tmp[2193]*kernel[4]+tmp[2194]*kernel[5]+tmp[2292]*kernel[6]+tmp[2293]*kernel[7]+tmp[2294]*kernel[8];
				ans[2194]<=tmp[2093]*kernel[0]+tmp[2094]*kernel[1]+tmp[2095]*kernel[2]+tmp[2193]*kernel[3]+tmp[2194]*kernel[4]+tmp[2195]*kernel[5]+tmp[2293]*kernel[6]+tmp[2294]*kernel[7]+tmp[2295]*kernel[8];
				ans[2195]<=tmp[2094]*kernel[0]+tmp[2095]*kernel[1]+tmp[2096]*kernel[2]+tmp[2194]*kernel[3]+tmp[2195]*kernel[4]+tmp[2196]*kernel[5]+tmp[2294]*kernel[6]+tmp[2295]*kernel[7]+tmp[2296]*kernel[8];
				ans[2196]<=tmp[2095]*kernel[0]+tmp[2096]*kernel[1]+tmp[2097]*kernel[2]+tmp[2195]*kernel[3]+tmp[2196]*kernel[4]+tmp[2197]*kernel[5]+tmp[2295]*kernel[6]+tmp[2296]*kernel[7]+tmp[2297]*kernel[8];
				ans[2197]<=tmp[2096]*kernel[0]+tmp[2097]*kernel[1]+tmp[2098]*kernel[2]+tmp[2196]*kernel[3]+tmp[2197]*kernel[4]+tmp[2198]*kernel[5]+tmp[2296]*kernel[6]+tmp[2297]*kernel[7]+tmp[2298]*kernel[8];
				ans[2198]<=tmp[2097]*kernel[0]+tmp[2098]*kernel[1]+tmp[2099]*kernel[2]+tmp[2197]*kernel[3]+tmp[2198]*kernel[4]+tmp[2199]*kernel[5]+tmp[2297]*kernel[6]+tmp[2298]*kernel[7]+tmp[2299]*kernel[8];
				ans[2199]<=tmp[2098]*kernel[0]+tmp[2099]*kernel[1]+tmp[2198]*kernel[3]+tmp[2199]*kernel[4]+tmp[2298]*kernel[6]+tmp[2299]*kernel[7];
				ans[2200]<=tmp[2100]*kernel[1]+tmp[2101]*kernel[2]+tmp[2200]*kernel[4]+tmp[2201]*kernel[5]+tmp[2300]*kernel[7]+tmp[2301]*kernel[8];
				ans[2201]<=tmp[2100]*kernel[0]+tmp[2101]*kernel[1]+tmp[2102]*kernel[2]+tmp[2200]*kernel[3]+tmp[2201]*kernel[4]+tmp[2202]*kernel[5]+tmp[2300]*kernel[6]+tmp[2301]*kernel[7]+tmp[2302]*kernel[8];
				ans[2202]<=tmp[2101]*kernel[0]+tmp[2102]*kernel[1]+tmp[2103]*kernel[2]+tmp[2201]*kernel[3]+tmp[2202]*kernel[4]+tmp[2203]*kernel[5]+tmp[2301]*kernel[6]+tmp[2302]*kernel[7]+tmp[2303]*kernel[8];
				ans[2203]<=tmp[2102]*kernel[0]+tmp[2103]*kernel[1]+tmp[2104]*kernel[2]+tmp[2202]*kernel[3]+tmp[2203]*kernel[4]+tmp[2204]*kernel[5]+tmp[2302]*kernel[6]+tmp[2303]*kernel[7]+tmp[2304]*kernel[8];
				ans[2204]<=tmp[2103]*kernel[0]+tmp[2104]*kernel[1]+tmp[2105]*kernel[2]+tmp[2203]*kernel[3]+tmp[2204]*kernel[4]+tmp[2205]*kernel[5]+tmp[2303]*kernel[6]+tmp[2304]*kernel[7]+tmp[2305]*kernel[8];
				ans[2205]<=tmp[2104]*kernel[0]+tmp[2105]*kernel[1]+tmp[2106]*kernel[2]+tmp[2204]*kernel[3]+tmp[2205]*kernel[4]+tmp[2206]*kernel[5]+tmp[2304]*kernel[6]+tmp[2305]*kernel[7]+tmp[2306]*kernel[8];
				ans[2206]<=tmp[2105]*kernel[0]+tmp[2106]*kernel[1]+tmp[2107]*kernel[2]+tmp[2205]*kernel[3]+tmp[2206]*kernel[4]+tmp[2207]*kernel[5]+tmp[2305]*kernel[6]+tmp[2306]*kernel[7]+tmp[2307]*kernel[8];
				ans[2207]<=tmp[2106]*kernel[0]+tmp[2107]*kernel[1]+tmp[2108]*kernel[2]+tmp[2206]*kernel[3]+tmp[2207]*kernel[4]+tmp[2208]*kernel[5]+tmp[2306]*kernel[6]+tmp[2307]*kernel[7]+tmp[2308]*kernel[8];
				ans[2208]<=tmp[2107]*kernel[0]+tmp[2108]*kernel[1]+tmp[2109]*kernel[2]+tmp[2207]*kernel[3]+tmp[2208]*kernel[4]+tmp[2209]*kernel[5]+tmp[2307]*kernel[6]+tmp[2308]*kernel[7]+tmp[2309]*kernel[8];
				ans[2209]<=tmp[2108]*kernel[0]+tmp[2109]*kernel[1]+tmp[2110]*kernel[2]+tmp[2208]*kernel[3]+tmp[2209]*kernel[4]+tmp[2210]*kernel[5]+tmp[2308]*kernel[6]+tmp[2309]*kernel[7]+tmp[2310]*kernel[8];
				ans[2210]<=tmp[2109]*kernel[0]+tmp[2110]*kernel[1]+tmp[2111]*kernel[2]+tmp[2209]*kernel[3]+tmp[2210]*kernel[4]+tmp[2211]*kernel[5]+tmp[2309]*kernel[6]+tmp[2310]*kernel[7]+tmp[2311]*kernel[8];
				ans[2211]<=tmp[2110]*kernel[0]+tmp[2111]*kernel[1]+tmp[2112]*kernel[2]+tmp[2210]*kernel[3]+tmp[2211]*kernel[4]+tmp[2212]*kernel[5]+tmp[2310]*kernel[6]+tmp[2311]*kernel[7]+tmp[2312]*kernel[8];
				ans[2212]<=tmp[2111]*kernel[0]+tmp[2112]*kernel[1]+tmp[2113]*kernel[2]+tmp[2211]*kernel[3]+tmp[2212]*kernel[4]+tmp[2213]*kernel[5]+tmp[2311]*kernel[6]+tmp[2312]*kernel[7]+tmp[2313]*kernel[8];
				ans[2213]<=tmp[2112]*kernel[0]+tmp[2113]*kernel[1]+tmp[2114]*kernel[2]+tmp[2212]*kernel[3]+tmp[2213]*kernel[4]+tmp[2214]*kernel[5]+tmp[2312]*kernel[6]+tmp[2313]*kernel[7]+tmp[2314]*kernel[8];
				ans[2214]<=tmp[2113]*kernel[0]+tmp[2114]*kernel[1]+tmp[2115]*kernel[2]+tmp[2213]*kernel[3]+tmp[2214]*kernel[4]+tmp[2215]*kernel[5]+tmp[2313]*kernel[6]+tmp[2314]*kernel[7]+tmp[2315]*kernel[8];
				ans[2215]<=tmp[2114]*kernel[0]+tmp[2115]*kernel[1]+tmp[2116]*kernel[2]+tmp[2214]*kernel[3]+tmp[2215]*kernel[4]+tmp[2216]*kernel[5]+tmp[2314]*kernel[6]+tmp[2315]*kernel[7]+tmp[2316]*kernel[8];
				ans[2216]<=tmp[2115]*kernel[0]+tmp[2116]*kernel[1]+tmp[2117]*kernel[2]+tmp[2215]*kernel[3]+tmp[2216]*kernel[4]+tmp[2217]*kernel[5]+tmp[2315]*kernel[6]+tmp[2316]*kernel[7]+tmp[2317]*kernel[8];
				ans[2217]<=tmp[2116]*kernel[0]+tmp[2117]*kernel[1]+tmp[2118]*kernel[2]+tmp[2216]*kernel[3]+tmp[2217]*kernel[4]+tmp[2218]*kernel[5]+tmp[2316]*kernel[6]+tmp[2317]*kernel[7]+tmp[2318]*kernel[8];
				ans[2218]<=tmp[2117]*kernel[0]+tmp[2118]*kernel[1]+tmp[2119]*kernel[2]+tmp[2217]*kernel[3]+tmp[2218]*kernel[4]+tmp[2219]*kernel[5]+tmp[2317]*kernel[6]+tmp[2318]*kernel[7]+tmp[2319]*kernel[8];
				ans[2219]<=tmp[2118]*kernel[0]+tmp[2119]*kernel[1]+tmp[2120]*kernel[2]+tmp[2218]*kernel[3]+tmp[2219]*kernel[4]+tmp[2220]*kernel[5]+tmp[2318]*kernel[6]+tmp[2319]*kernel[7]+tmp[2320]*kernel[8];
				ans[2220]<=tmp[2119]*kernel[0]+tmp[2120]*kernel[1]+tmp[2121]*kernel[2]+tmp[2219]*kernel[3]+tmp[2220]*kernel[4]+tmp[2221]*kernel[5]+tmp[2319]*kernel[6]+tmp[2320]*kernel[7]+tmp[2321]*kernel[8];
				ans[2221]<=tmp[2120]*kernel[0]+tmp[2121]*kernel[1]+tmp[2122]*kernel[2]+tmp[2220]*kernel[3]+tmp[2221]*kernel[4]+tmp[2222]*kernel[5]+tmp[2320]*kernel[6]+tmp[2321]*kernel[7]+tmp[2322]*kernel[8];
				ans[2222]<=tmp[2121]*kernel[0]+tmp[2122]*kernel[1]+tmp[2123]*kernel[2]+tmp[2221]*kernel[3]+tmp[2222]*kernel[4]+tmp[2223]*kernel[5]+tmp[2321]*kernel[6]+tmp[2322]*kernel[7]+tmp[2323]*kernel[8];
				ans[2223]<=tmp[2122]*kernel[0]+tmp[2123]*kernel[1]+tmp[2124]*kernel[2]+tmp[2222]*kernel[3]+tmp[2223]*kernel[4]+tmp[2224]*kernel[5]+tmp[2322]*kernel[6]+tmp[2323]*kernel[7]+tmp[2324]*kernel[8];
				ans[2224]<=tmp[2123]*kernel[0]+tmp[2124]*kernel[1]+tmp[2125]*kernel[2]+tmp[2223]*kernel[3]+tmp[2224]*kernel[4]+tmp[2225]*kernel[5]+tmp[2323]*kernel[6]+tmp[2324]*kernel[7]+tmp[2325]*kernel[8];
				ans[2225]<=tmp[2124]*kernel[0]+tmp[2125]*kernel[1]+tmp[2126]*kernel[2]+tmp[2224]*kernel[3]+tmp[2225]*kernel[4]+tmp[2226]*kernel[5]+tmp[2324]*kernel[6]+tmp[2325]*kernel[7]+tmp[2326]*kernel[8];
				ans[2226]<=tmp[2125]*kernel[0]+tmp[2126]*kernel[1]+tmp[2127]*kernel[2]+tmp[2225]*kernel[3]+tmp[2226]*kernel[4]+tmp[2227]*kernel[5]+tmp[2325]*kernel[6]+tmp[2326]*kernel[7]+tmp[2327]*kernel[8];
				ans[2227]<=tmp[2126]*kernel[0]+tmp[2127]*kernel[1]+tmp[2128]*kernel[2]+tmp[2226]*kernel[3]+tmp[2227]*kernel[4]+tmp[2228]*kernel[5]+tmp[2326]*kernel[6]+tmp[2327]*kernel[7]+tmp[2328]*kernel[8];
				ans[2228]<=tmp[2127]*kernel[0]+tmp[2128]*kernel[1]+tmp[2129]*kernel[2]+tmp[2227]*kernel[3]+tmp[2228]*kernel[4]+tmp[2229]*kernel[5]+tmp[2327]*kernel[6]+tmp[2328]*kernel[7]+tmp[2329]*kernel[8];
				ans[2229]<=tmp[2128]*kernel[0]+tmp[2129]*kernel[1]+tmp[2130]*kernel[2]+tmp[2228]*kernel[3]+tmp[2229]*kernel[4]+tmp[2230]*kernel[5]+tmp[2328]*kernel[6]+tmp[2329]*kernel[7]+tmp[2330]*kernel[8];
				ans[2230]<=tmp[2129]*kernel[0]+tmp[2130]*kernel[1]+tmp[2131]*kernel[2]+tmp[2229]*kernel[3]+tmp[2230]*kernel[4]+tmp[2231]*kernel[5]+tmp[2329]*kernel[6]+tmp[2330]*kernel[7]+tmp[2331]*kernel[8];
				ans[2231]<=tmp[2130]*kernel[0]+tmp[2131]*kernel[1]+tmp[2132]*kernel[2]+tmp[2230]*kernel[3]+tmp[2231]*kernel[4]+tmp[2232]*kernel[5]+tmp[2330]*kernel[6]+tmp[2331]*kernel[7]+tmp[2332]*kernel[8];
				ans[2232]<=tmp[2131]*kernel[0]+tmp[2132]*kernel[1]+tmp[2133]*kernel[2]+tmp[2231]*kernel[3]+tmp[2232]*kernel[4]+tmp[2233]*kernel[5]+tmp[2331]*kernel[6]+tmp[2332]*kernel[7]+tmp[2333]*kernel[8];
				ans[2233]<=tmp[2132]*kernel[0]+tmp[2133]*kernel[1]+tmp[2134]*kernel[2]+tmp[2232]*kernel[3]+tmp[2233]*kernel[4]+tmp[2234]*kernel[5]+tmp[2332]*kernel[6]+tmp[2333]*kernel[7]+tmp[2334]*kernel[8];
				ans[2234]<=tmp[2133]*kernel[0]+tmp[2134]*kernel[1]+tmp[2135]*kernel[2]+tmp[2233]*kernel[3]+tmp[2234]*kernel[4]+tmp[2235]*kernel[5]+tmp[2333]*kernel[6]+tmp[2334]*kernel[7]+tmp[2335]*kernel[8];
				ans[2235]<=tmp[2134]*kernel[0]+tmp[2135]*kernel[1]+tmp[2136]*kernel[2]+tmp[2234]*kernel[3]+tmp[2235]*kernel[4]+tmp[2236]*kernel[5]+tmp[2334]*kernel[6]+tmp[2335]*kernel[7]+tmp[2336]*kernel[8];
				ans[2236]<=tmp[2135]*kernel[0]+tmp[2136]*kernel[1]+tmp[2137]*kernel[2]+tmp[2235]*kernel[3]+tmp[2236]*kernel[4]+tmp[2237]*kernel[5]+tmp[2335]*kernel[6]+tmp[2336]*kernel[7]+tmp[2337]*kernel[8];
				ans[2237]<=tmp[2136]*kernel[0]+tmp[2137]*kernel[1]+tmp[2138]*kernel[2]+tmp[2236]*kernel[3]+tmp[2237]*kernel[4]+tmp[2238]*kernel[5]+tmp[2336]*kernel[6]+tmp[2337]*kernel[7]+tmp[2338]*kernel[8];
				ans[2238]<=tmp[2137]*kernel[0]+tmp[2138]*kernel[1]+tmp[2139]*kernel[2]+tmp[2237]*kernel[3]+tmp[2238]*kernel[4]+tmp[2239]*kernel[5]+tmp[2337]*kernel[6]+tmp[2338]*kernel[7]+tmp[2339]*kernel[8];
				ans[2239]<=tmp[2138]*kernel[0]+tmp[2139]*kernel[1]+tmp[2140]*kernel[2]+tmp[2238]*kernel[3]+tmp[2239]*kernel[4]+tmp[2240]*kernel[5]+tmp[2338]*kernel[6]+tmp[2339]*kernel[7]+tmp[2340]*kernel[8];
				ans[2240]<=tmp[2139]*kernel[0]+tmp[2140]*kernel[1]+tmp[2141]*kernel[2]+tmp[2239]*kernel[3]+tmp[2240]*kernel[4]+tmp[2241]*kernel[5]+tmp[2339]*kernel[6]+tmp[2340]*kernel[7]+tmp[2341]*kernel[8];
				ans[2241]<=tmp[2140]*kernel[0]+tmp[2141]*kernel[1]+tmp[2142]*kernel[2]+tmp[2240]*kernel[3]+tmp[2241]*kernel[4]+tmp[2242]*kernel[5]+tmp[2340]*kernel[6]+tmp[2341]*kernel[7]+tmp[2342]*kernel[8];
				ans[2242]<=tmp[2141]*kernel[0]+tmp[2142]*kernel[1]+tmp[2143]*kernel[2]+tmp[2241]*kernel[3]+tmp[2242]*kernel[4]+tmp[2243]*kernel[5]+tmp[2341]*kernel[6]+tmp[2342]*kernel[7]+tmp[2343]*kernel[8];
				ans[2243]<=tmp[2142]*kernel[0]+tmp[2143]*kernel[1]+tmp[2144]*kernel[2]+tmp[2242]*kernel[3]+tmp[2243]*kernel[4]+tmp[2244]*kernel[5]+tmp[2342]*kernel[6]+tmp[2343]*kernel[7]+tmp[2344]*kernel[8];
				ans[2244]<=tmp[2143]*kernel[0]+tmp[2144]*kernel[1]+tmp[2145]*kernel[2]+tmp[2243]*kernel[3]+tmp[2244]*kernel[4]+tmp[2245]*kernel[5]+tmp[2343]*kernel[6]+tmp[2344]*kernel[7]+tmp[2345]*kernel[8];
				ans[2245]<=tmp[2144]*kernel[0]+tmp[2145]*kernel[1]+tmp[2146]*kernel[2]+tmp[2244]*kernel[3]+tmp[2245]*kernel[4]+tmp[2246]*kernel[5]+tmp[2344]*kernel[6]+tmp[2345]*kernel[7]+tmp[2346]*kernel[8];
				ans[2246]<=tmp[2145]*kernel[0]+tmp[2146]*kernel[1]+tmp[2147]*kernel[2]+tmp[2245]*kernel[3]+tmp[2246]*kernel[4]+tmp[2247]*kernel[5]+tmp[2345]*kernel[6]+tmp[2346]*kernel[7]+tmp[2347]*kernel[8];
				ans[2247]<=tmp[2146]*kernel[0]+tmp[2147]*kernel[1]+tmp[2148]*kernel[2]+tmp[2246]*kernel[3]+tmp[2247]*kernel[4]+tmp[2248]*kernel[5]+tmp[2346]*kernel[6]+tmp[2347]*kernel[7]+tmp[2348]*kernel[8];
				ans[2248]<=tmp[2147]*kernel[0]+tmp[2148]*kernel[1]+tmp[2149]*kernel[2]+tmp[2247]*kernel[3]+tmp[2248]*kernel[4]+tmp[2249]*kernel[5]+tmp[2347]*kernel[6]+tmp[2348]*kernel[7]+tmp[2349]*kernel[8];
				ans[2249]<=tmp[2148]*kernel[0]+tmp[2149]*kernel[1]+tmp[2150]*kernel[2]+tmp[2248]*kernel[3]+tmp[2249]*kernel[4]+tmp[2250]*kernel[5]+tmp[2348]*kernel[6]+tmp[2349]*kernel[7]+tmp[2350]*kernel[8];
				ans[2250]<=tmp[2149]*kernel[0]+tmp[2150]*kernel[1]+tmp[2151]*kernel[2]+tmp[2249]*kernel[3]+tmp[2250]*kernel[4]+tmp[2251]*kernel[5]+tmp[2349]*kernel[6]+tmp[2350]*kernel[7]+tmp[2351]*kernel[8];
				ans[2251]<=tmp[2150]*kernel[0]+tmp[2151]*kernel[1]+tmp[2152]*kernel[2]+tmp[2250]*kernel[3]+tmp[2251]*kernel[4]+tmp[2252]*kernel[5]+tmp[2350]*kernel[6]+tmp[2351]*kernel[7]+tmp[2352]*kernel[8];
				ans[2252]<=tmp[2151]*kernel[0]+tmp[2152]*kernel[1]+tmp[2153]*kernel[2]+tmp[2251]*kernel[3]+tmp[2252]*kernel[4]+tmp[2253]*kernel[5]+tmp[2351]*kernel[6]+tmp[2352]*kernel[7]+tmp[2353]*kernel[8];
				ans[2253]<=tmp[2152]*kernel[0]+tmp[2153]*kernel[1]+tmp[2154]*kernel[2]+tmp[2252]*kernel[3]+tmp[2253]*kernel[4]+tmp[2254]*kernel[5]+tmp[2352]*kernel[6]+tmp[2353]*kernel[7]+tmp[2354]*kernel[8];
				ans[2254]<=tmp[2153]*kernel[0]+tmp[2154]*kernel[1]+tmp[2155]*kernel[2]+tmp[2253]*kernel[3]+tmp[2254]*kernel[4]+tmp[2255]*kernel[5]+tmp[2353]*kernel[6]+tmp[2354]*kernel[7]+tmp[2355]*kernel[8];
				ans[2255]<=tmp[2154]*kernel[0]+tmp[2155]*kernel[1]+tmp[2156]*kernel[2]+tmp[2254]*kernel[3]+tmp[2255]*kernel[4]+tmp[2256]*kernel[5]+tmp[2354]*kernel[6]+tmp[2355]*kernel[7]+tmp[2356]*kernel[8];
				ans[2256]<=tmp[2155]*kernel[0]+tmp[2156]*kernel[1]+tmp[2157]*kernel[2]+tmp[2255]*kernel[3]+tmp[2256]*kernel[4]+tmp[2257]*kernel[5]+tmp[2355]*kernel[6]+tmp[2356]*kernel[7]+tmp[2357]*kernel[8];
				ans[2257]<=tmp[2156]*kernel[0]+tmp[2157]*kernel[1]+tmp[2158]*kernel[2]+tmp[2256]*kernel[3]+tmp[2257]*kernel[4]+tmp[2258]*kernel[5]+tmp[2356]*kernel[6]+tmp[2357]*kernel[7]+tmp[2358]*kernel[8];
				ans[2258]<=tmp[2157]*kernel[0]+tmp[2158]*kernel[1]+tmp[2159]*kernel[2]+tmp[2257]*kernel[3]+tmp[2258]*kernel[4]+tmp[2259]*kernel[5]+tmp[2357]*kernel[6]+tmp[2358]*kernel[7]+tmp[2359]*kernel[8];
				ans[2259]<=tmp[2158]*kernel[0]+tmp[2159]*kernel[1]+tmp[2160]*kernel[2]+tmp[2258]*kernel[3]+tmp[2259]*kernel[4]+tmp[2260]*kernel[5]+tmp[2358]*kernel[6]+tmp[2359]*kernel[7]+tmp[2360]*kernel[8];
				ans[2260]<=tmp[2159]*kernel[0]+tmp[2160]*kernel[1]+tmp[2161]*kernel[2]+tmp[2259]*kernel[3]+tmp[2260]*kernel[4]+tmp[2261]*kernel[5]+tmp[2359]*kernel[6]+tmp[2360]*kernel[7]+tmp[2361]*kernel[8];
				ans[2261]<=tmp[2160]*kernel[0]+tmp[2161]*kernel[1]+tmp[2162]*kernel[2]+tmp[2260]*kernel[3]+tmp[2261]*kernel[4]+tmp[2262]*kernel[5]+tmp[2360]*kernel[6]+tmp[2361]*kernel[7]+tmp[2362]*kernel[8];
				ans[2262]<=tmp[2161]*kernel[0]+tmp[2162]*kernel[1]+tmp[2163]*kernel[2]+tmp[2261]*kernel[3]+tmp[2262]*kernel[4]+tmp[2263]*kernel[5]+tmp[2361]*kernel[6]+tmp[2362]*kernel[7]+tmp[2363]*kernel[8];
				ans[2263]<=tmp[2162]*kernel[0]+tmp[2163]*kernel[1]+tmp[2164]*kernel[2]+tmp[2262]*kernel[3]+tmp[2263]*kernel[4]+tmp[2264]*kernel[5]+tmp[2362]*kernel[6]+tmp[2363]*kernel[7]+tmp[2364]*kernel[8];
				ans[2264]<=tmp[2163]*kernel[0]+tmp[2164]*kernel[1]+tmp[2165]*kernel[2]+tmp[2263]*kernel[3]+tmp[2264]*kernel[4]+tmp[2265]*kernel[5]+tmp[2363]*kernel[6]+tmp[2364]*kernel[7]+tmp[2365]*kernel[8];
				ans[2265]<=tmp[2164]*kernel[0]+tmp[2165]*kernel[1]+tmp[2166]*kernel[2]+tmp[2264]*kernel[3]+tmp[2265]*kernel[4]+tmp[2266]*kernel[5]+tmp[2364]*kernel[6]+tmp[2365]*kernel[7]+tmp[2366]*kernel[8];
				ans[2266]<=tmp[2165]*kernel[0]+tmp[2166]*kernel[1]+tmp[2167]*kernel[2]+tmp[2265]*kernel[3]+tmp[2266]*kernel[4]+tmp[2267]*kernel[5]+tmp[2365]*kernel[6]+tmp[2366]*kernel[7]+tmp[2367]*kernel[8];
				ans[2267]<=tmp[2166]*kernel[0]+tmp[2167]*kernel[1]+tmp[2168]*kernel[2]+tmp[2266]*kernel[3]+tmp[2267]*kernel[4]+tmp[2268]*kernel[5]+tmp[2366]*kernel[6]+tmp[2367]*kernel[7]+tmp[2368]*kernel[8];
				ans[2268]<=tmp[2167]*kernel[0]+tmp[2168]*kernel[1]+tmp[2169]*kernel[2]+tmp[2267]*kernel[3]+tmp[2268]*kernel[4]+tmp[2269]*kernel[5]+tmp[2367]*kernel[6]+tmp[2368]*kernel[7]+tmp[2369]*kernel[8];
				ans[2269]<=tmp[2168]*kernel[0]+tmp[2169]*kernel[1]+tmp[2170]*kernel[2]+tmp[2268]*kernel[3]+tmp[2269]*kernel[4]+tmp[2270]*kernel[5]+tmp[2368]*kernel[6]+tmp[2369]*kernel[7]+tmp[2370]*kernel[8];
				ans[2270]<=tmp[2169]*kernel[0]+tmp[2170]*kernel[1]+tmp[2171]*kernel[2]+tmp[2269]*kernel[3]+tmp[2270]*kernel[4]+tmp[2271]*kernel[5]+tmp[2369]*kernel[6]+tmp[2370]*kernel[7]+tmp[2371]*kernel[8];
				ans[2271]<=tmp[2170]*kernel[0]+tmp[2171]*kernel[1]+tmp[2172]*kernel[2]+tmp[2270]*kernel[3]+tmp[2271]*kernel[4]+tmp[2272]*kernel[5]+tmp[2370]*kernel[6]+tmp[2371]*kernel[7]+tmp[2372]*kernel[8];
				ans[2272]<=tmp[2171]*kernel[0]+tmp[2172]*kernel[1]+tmp[2173]*kernel[2]+tmp[2271]*kernel[3]+tmp[2272]*kernel[4]+tmp[2273]*kernel[5]+tmp[2371]*kernel[6]+tmp[2372]*kernel[7]+tmp[2373]*kernel[8];
				ans[2273]<=tmp[2172]*kernel[0]+tmp[2173]*kernel[1]+tmp[2174]*kernel[2]+tmp[2272]*kernel[3]+tmp[2273]*kernel[4]+tmp[2274]*kernel[5]+tmp[2372]*kernel[6]+tmp[2373]*kernel[7]+tmp[2374]*kernel[8];
				ans[2274]<=tmp[2173]*kernel[0]+tmp[2174]*kernel[1]+tmp[2175]*kernel[2]+tmp[2273]*kernel[3]+tmp[2274]*kernel[4]+tmp[2275]*kernel[5]+tmp[2373]*kernel[6]+tmp[2374]*kernel[7]+tmp[2375]*kernel[8];
				ans[2275]<=tmp[2174]*kernel[0]+tmp[2175]*kernel[1]+tmp[2176]*kernel[2]+tmp[2274]*kernel[3]+tmp[2275]*kernel[4]+tmp[2276]*kernel[5]+tmp[2374]*kernel[6]+tmp[2375]*kernel[7]+tmp[2376]*kernel[8];
				ans[2276]<=tmp[2175]*kernel[0]+tmp[2176]*kernel[1]+tmp[2177]*kernel[2]+tmp[2275]*kernel[3]+tmp[2276]*kernel[4]+tmp[2277]*kernel[5]+tmp[2375]*kernel[6]+tmp[2376]*kernel[7]+tmp[2377]*kernel[8];
				ans[2277]<=tmp[2176]*kernel[0]+tmp[2177]*kernel[1]+tmp[2178]*kernel[2]+tmp[2276]*kernel[3]+tmp[2277]*kernel[4]+tmp[2278]*kernel[5]+tmp[2376]*kernel[6]+tmp[2377]*kernel[7]+tmp[2378]*kernel[8];
				ans[2278]<=tmp[2177]*kernel[0]+tmp[2178]*kernel[1]+tmp[2179]*kernel[2]+tmp[2277]*kernel[3]+tmp[2278]*kernel[4]+tmp[2279]*kernel[5]+tmp[2377]*kernel[6]+tmp[2378]*kernel[7]+tmp[2379]*kernel[8];
				ans[2279]<=tmp[2178]*kernel[0]+tmp[2179]*kernel[1]+tmp[2180]*kernel[2]+tmp[2278]*kernel[3]+tmp[2279]*kernel[4]+tmp[2280]*kernel[5]+tmp[2378]*kernel[6]+tmp[2379]*kernel[7]+tmp[2380]*kernel[8];
				ans[2280]<=tmp[2179]*kernel[0]+tmp[2180]*kernel[1]+tmp[2181]*kernel[2]+tmp[2279]*kernel[3]+tmp[2280]*kernel[4]+tmp[2281]*kernel[5]+tmp[2379]*kernel[6]+tmp[2380]*kernel[7]+tmp[2381]*kernel[8];
				ans[2281]<=tmp[2180]*kernel[0]+tmp[2181]*kernel[1]+tmp[2182]*kernel[2]+tmp[2280]*kernel[3]+tmp[2281]*kernel[4]+tmp[2282]*kernel[5]+tmp[2380]*kernel[6]+tmp[2381]*kernel[7]+tmp[2382]*kernel[8];
				ans[2282]<=tmp[2181]*kernel[0]+tmp[2182]*kernel[1]+tmp[2183]*kernel[2]+tmp[2281]*kernel[3]+tmp[2282]*kernel[4]+tmp[2283]*kernel[5]+tmp[2381]*kernel[6]+tmp[2382]*kernel[7]+tmp[2383]*kernel[8];
				ans[2283]<=tmp[2182]*kernel[0]+tmp[2183]*kernel[1]+tmp[2184]*kernel[2]+tmp[2282]*kernel[3]+tmp[2283]*kernel[4]+tmp[2284]*kernel[5]+tmp[2382]*kernel[6]+tmp[2383]*kernel[7]+tmp[2384]*kernel[8];
				ans[2284]<=tmp[2183]*kernel[0]+tmp[2184]*kernel[1]+tmp[2185]*kernel[2]+tmp[2283]*kernel[3]+tmp[2284]*kernel[4]+tmp[2285]*kernel[5]+tmp[2383]*kernel[6]+tmp[2384]*kernel[7]+tmp[2385]*kernel[8];
				ans[2285]<=tmp[2184]*kernel[0]+tmp[2185]*kernel[1]+tmp[2186]*kernel[2]+tmp[2284]*kernel[3]+tmp[2285]*kernel[4]+tmp[2286]*kernel[5]+tmp[2384]*kernel[6]+tmp[2385]*kernel[7]+tmp[2386]*kernel[8];
				ans[2286]<=tmp[2185]*kernel[0]+tmp[2186]*kernel[1]+tmp[2187]*kernel[2]+tmp[2285]*kernel[3]+tmp[2286]*kernel[4]+tmp[2287]*kernel[5]+tmp[2385]*kernel[6]+tmp[2386]*kernel[7]+tmp[2387]*kernel[8];
				ans[2287]<=tmp[2186]*kernel[0]+tmp[2187]*kernel[1]+tmp[2188]*kernel[2]+tmp[2286]*kernel[3]+tmp[2287]*kernel[4]+tmp[2288]*kernel[5]+tmp[2386]*kernel[6]+tmp[2387]*kernel[7]+tmp[2388]*kernel[8];
				ans[2288]<=tmp[2187]*kernel[0]+tmp[2188]*kernel[1]+tmp[2189]*kernel[2]+tmp[2287]*kernel[3]+tmp[2288]*kernel[4]+tmp[2289]*kernel[5]+tmp[2387]*kernel[6]+tmp[2388]*kernel[7]+tmp[2389]*kernel[8];
				ans[2289]<=tmp[2188]*kernel[0]+tmp[2189]*kernel[1]+tmp[2190]*kernel[2]+tmp[2288]*kernel[3]+tmp[2289]*kernel[4]+tmp[2290]*kernel[5]+tmp[2388]*kernel[6]+tmp[2389]*kernel[7]+tmp[2390]*kernel[8];
				ans[2290]<=tmp[2189]*kernel[0]+tmp[2190]*kernel[1]+tmp[2191]*kernel[2]+tmp[2289]*kernel[3]+tmp[2290]*kernel[4]+tmp[2291]*kernel[5]+tmp[2389]*kernel[6]+tmp[2390]*kernel[7]+tmp[2391]*kernel[8];
				ans[2291]<=tmp[2190]*kernel[0]+tmp[2191]*kernel[1]+tmp[2192]*kernel[2]+tmp[2290]*kernel[3]+tmp[2291]*kernel[4]+tmp[2292]*kernel[5]+tmp[2390]*kernel[6]+tmp[2391]*kernel[7]+tmp[2392]*kernel[8];
				ans[2292]<=tmp[2191]*kernel[0]+tmp[2192]*kernel[1]+tmp[2193]*kernel[2]+tmp[2291]*kernel[3]+tmp[2292]*kernel[4]+tmp[2293]*kernel[5]+tmp[2391]*kernel[6]+tmp[2392]*kernel[7]+tmp[2393]*kernel[8];
				ans[2293]<=tmp[2192]*kernel[0]+tmp[2193]*kernel[1]+tmp[2194]*kernel[2]+tmp[2292]*kernel[3]+tmp[2293]*kernel[4]+tmp[2294]*kernel[5]+tmp[2392]*kernel[6]+tmp[2393]*kernel[7]+tmp[2394]*kernel[8];
				ans[2294]<=tmp[2193]*kernel[0]+tmp[2194]*kernel[1]+tmp[2195]*kernel[2]+tmp[2293]*kernel[3]+tmp[2294]*kernel[4]+tmp[2295]*kernel[5]+tmp[2393]*kernel[6]+tmp[2394]*kernel[7]+tmp[2395]*kernel[8];
				ans[2295]<=tmp[2194]*kernel[0]+tmp[2195]*kernel[1]+tmp[2196]*kernel[2]+tmp[2294]*kernel[3]+tmp[2295]*kernel[4]+tmp[2296]*kernel[5]+tmp[2394]*kernel[6]+tmp[2395]*kernel[7]+tmp[2396]*kernel[8];
				ans[2296]<=tmp[2195]*kernel[0]+tmp[2196]*kernel[1]+tmp[2197]*kernel[2]+tmp[2295]*kernel[3]+tmp[2296]*kernel[4]+tmp[2297]*kernel[5]+tmp[2395]*kernel[6]+tmp[2396]*kernel[7]+tmp[2397]*kernel[8];
				ans[2297]<=tmp[2196]*kernel[0]+tmp[2197]*kernel[1]+tmp[2198]*kernel[2]+tmp[2296]*kernel[3]+tmp[2297]*kernel[4]+tmp[2298]*kernel[5]+tmp[2396]*kernel[6]+tmp[2397]*kernel[7]+tmp[2398]*kernel[8];
				ans[2298]<=tmp[2197]*kernel[0]+tmp[2198]*kernel[1]+tmp[2199]*kernel[2]+tmp[2297]*kernel[3]+tmp[2298]*kernel[4]+tmp[2299]*kernel[5]+tmp[2397]*kernel[6]+tmp[2398]*kernel[7]+tmp[2399]*kernel[8];
				ans[2299]<=tmp[2198]*kernel[0]+tmp[2199]*kernel[1]+tmp[2298]*kernel[3]+tmp[2299]*kernel[4]+tmp[2398]*kernel[6]+tmp[2399]*kernel[7];
				ans[2300]<=tmp[2200]*kernel[1]+tmp[2201]*kernel[2]+tmp[2300]*kernel[4]+tmp[2301]*kernel[5]+tmp[2400]*kernel[7]+tmp[2401]*kernel[8];
				ans[2301]<=tmp[2200]*kernel[0]+tmp[2201]*kernel[1]+tmp[2202]*kernel[2]+tmp[2300]*kernel[3]+tmp[2301]*kernel[4]+tmp[2302]*kernel[5]+tmp[2400]*kernel[6]+tmp[2401]*kernel[7]+tmp[2402]*kernel[8];
				ans[2302]<=tmp[2201]*kernel[0]+tmp[2202]*kernel[1]+tmp[2203]*kernel[2]+tmp[2301]*kernel[3]+tmp[2302]*kernel[4]+tmp[2303]*kernel[5]+tmp[2401]*kernel[6]+tmp[2402]*kernel[7]+tmp[2403]*kernel[8];
				ans[2303]<=tmp[2202]*kernel[0]+tmp[2203]*kernel[1]+tmp[2204]*kernel[2]+tmp[2302]*kernel[3]+tmp[2303]*kernel[4]+tmp[2304]*kernel[5]+tmp[2402]*kernel[6]+tmp[2403]*kernel[7]+tmp[2404]*kernel[8];
				ans[2304]<=tmp[2203]*kernel[0]+tmp[2204]*kernel[1]+tmp[2205]*kernel[2]+tmp[2303]*kernel[3]+tmp[2304]*kernel[4]+tmp[2305]*kernel[5]+tmp[2403]*kernel[6]+tmp[2404]*kernel[7]+tmp[2405]*kernel[8];
				ans[2305]<=tmp[2204]*kernel[0]+tmp[2205]*kernel[1]+tmp[2206]*kernel[2]+tmp[2304]*kernel[3]+tmp[2305]*kernel[4]+tmp[2306]*kernel[5]+tmp[2404]*kernel[6]+tmp[2405]*kernel[7]+tmp[2406]*kernel[8];
				ans[2306]<=tmp[2205]*kernel[0]+tmp[2206]*kernel[1]+tmp[2207]*kernel[2]+tmp[2305]*kernel[3]+tmp[2306]*kernel[4]+tmp[2307]*kernel[5]+tmp[2405]*kernel[6]+tmp[2406]*kernel[7]+tmp[2407]*kernel[8];
				ans[2307]<=tmp[2206]*kernel[0]+tmp[2207]*kernel[1]+tmp[2208]*kernel[2]+tmp[2306]*kernel[3]+tmp[2307]*kernel[4]+tmp[2308]*kernel[5]+tmp[2406]*kernel[6]+tmp[2407]*kernel[7]+tmp[2408]*kernel[8];
				ans[2308]<=tmp[2207]*kernel[0]+tmp[2208]*kernel[1]+tmp[2209]*kernel[2]+tmp[2307]*kernel[3]+tmp[2308]*kernel[4]+tmp[2309]*kernel[5]+tmp[2407]*kernel[6]+tmp[2408]*kernel[7]+tmp[2409]*kernel[8];
				ans[2309]<=tmp[2208]*kernel[0]+tmp[2209]*kernel[1]+tmp[2210]*kernel[2]+tmp[2308]*kernel[3]+tmp[2309]*kernel[4]+tmp[2310]*kernel[5]+tmp[2408]*kernel[6]+tmp[2409]*kernel[7]+tmp[2410]*kernel[8];
				ans[2310]<=tmp[2209]*kernel[0]+tmp[2210]*kernel[1]+tmp[2211]*kernel[2]+tmp[2309]*kernel[3]+tmp[2310]*kernel[4]+tmp[2311]*kernel[5]+tmp[2409]*kernel[6]+tmp[2410]*kernel[7]+tmp[2411]*kernel[8];
				ans[2311]<=tmp[2210]*kernel[0]+tmp[2211]*kernel[1]+tmp[2212]*kernel[2]+tmp[2310]*kernel[3]+tmp[2311]*kernel[4]+tmp[2312]*kernel[5]+tmp[2410]*kernel[6]+tmp[2411]*kernel[7]+tmp[2412]*kernel[8];
				ans[2312]<=tmp[2211]*kernel[0]+tmp[2212]*kernel[1]+tmp[2213]*kernel[2]+tmp[2311]*kernel[3]+tmp[2312]*kernel[4]+tmp[2313]*kernel[5]+tmp[2411]*kernel[6]+tmp[2412]*kernel[7]+tmp[2413]*kernel[8];
				ans[2313]<=tmp[2212]*kernel[0]+tmp[2213]*kernel[1]+tmp[2214]*kernel[2]+tmp[2312]*kernel[3]+tmp[2313]*kernel[4]+tmp[2314]*kernel[5]+tmp[2412]*kernel[6]+tmp[2413]*kernel[7]+tmp[2414]*kernel[8];
				ans[2314]<=tmp[2213]*kernel[0]+tmp[2214]*kernel[1]+tmp[2215]*kernel[2]+tmp[2313]*kernel[3]+tmp[2314]*kernel[4]+tmp[2315]*kernel[5]+tmp[2413]*kernel[6]+tmp[2414]*kernel[7]+tmp[2415]*kernel[8];
				ans[2315]<=tmp[2214]*kernel[0]+tmp[2215]*kernel[1]+tmp[2216]*kernel[2]+tmp[2314]*kernel[3]+tmp[2315]*kernel[4]+tmp[2316]*kernel[5]+tmp[2414]*kernel[6]+tmp[2415]*kernel[7]+tmp[2416]*kernel[8];
				ans[2316]<=tmp[2215]*kernel[0]+tmp[2216]*kernel[1]+tmp[2217]*kernel[2]+tmp[2315]*kernel[3]+tmp[2316]*kernel[4]+tmp[2317]*kernel[5]+tmp[2415]*kernel[6]+tmp[2416]*kernel[7]+tmp[2417]*kernel[8];
				ans[2317]<=tmp[2216]*kernel[0]+tmp[2217]*kernel[1]+tmp[2218]*kernel[2]+tmp[2316]*kernel[3]+tmp[2317]*kernel[4]+tmp[2318]*kernel[5]+tmp[2416]*kernel[6]+tmp[2417]*kernel[7]+tmp[2418]*kernel[8];
				ans[2318]<=tmp[2217]*kernel[0]+tmp[2218]*kernel[1]+tmp[2219]*kernel[2]+tmp[2317]*kernel[3]+tmp[2318]*kernel[4]+tmp[2319]*kernel[5]+tmp[2417]*kernel[6]+tmp[2418]*kernel[7]+tmp[2419]*kernel[8];
				ans[2319]<=tmp[2218]*kernel[0]+tmp[2219]*kernel[1]+tmp[2220]*kernel[2]+tmp[2318]*kernel[3]+tmp[2319]*kernel[4]+tmp[2320]*kernel[5]+tmp[2418]*kernel[6]+tmp[2419]*kernel[7]+tmp[2420]*kernel[8];
				ans[2320]<=tmp[2219]*kernel[0]+tmp[2220]*kernel[1]+tmp[2221]*kernel[2]+tmp[2319]*kernel[3]+tmp[2320]*kernel[4]+tmp[2321]*kernel[5]+tmp[2419]*kernel[6]+tmp[2420]*kernel[7]+tmp[2421]*kernel[8];
				ans[2321]<=tmp[2220]*kernel[0]+tmp[2221]*kernel[1]+tmp[2222]*kernel[2]+tmp[2320]*kernel[3]+tmp[2321]*kernel[4]+tmp[2322]*kernel[5]+tmp[2420]*kernel[6]+tmp[2421]*kernel[7]+tmp[2422]*kernel[8];
				ans[2322]<=tmp[2221]*kernel[0]+tmp[2222]*kernel[1]+tmp[2223]*kernel[2]+tmp[2321]*kernel[3]+tmp[2322]*kernel[4]+tmp[2323]*kernel[5]+tmp[2421]*kernel[6]+tmp[2422]*kernel[7]+tmp[2423]*kernel[8];
				ans[2323]<=tmp[2222]*kernel[0]+tmp[2223]*kernel[1]+tmp[2224]*kernel[2]+tmp[2322]*kernel[3]+tmp[2323]*kernel[4]+tmp[2324]*kernel[5]+tmp[2422]*kernel[6]+tmp[2423]*kernel[7]+tmp[2424]*kernel[8];
				ans[2324]<=tmp[2223]*kernel[0]+tmp[2224]*kernel[1]+tmp[2225]*kernel[2]+tmp[2323]*kernel[3]+tmp[2324]*kernel[4]+tmp[2325]*kernel[5]+tmp[2423]*kernel[6]+tmp[2424]*kernel[7]+tmp[2425]*kernel[8];
				ans[2325]<=tmp[2224]*kernel[0]+tmp[2225]*kernel[1]+tmp[2226]*kernel[2]+tmp[2324]*kernel[3]+tmp[2325]*kernel[4]+tmp[2326]*kernel[5]+tmp[2424]*kernel[6]+tmp[2425]*kernel[7]+tmp[2426]*kernel[8];
				ans[2326]<=tmp[2225]*kernel[0]+tmp[2226]*kernel[1]+tmp[2227]*kernel[2]+tmp[2325]*kernel[3]+tmp[2326]*kernel[4]+tmp[2327]*kernel[5]+tmp[2425]*kernel[6]+tmp[2426]*kernel[7]+tmp[2427]*kernel[8];
				ans[2327]<=tmp[2226]*kernel[0]+tmp[2227]*kernel[1]+tmp[2228]*kernel[2]+tmp[2326]*kernel[3]+tmp[2327]*kernel[4]+tmp[2328]*kernel[5]+tmp[2426]*kernel[6]+tmp[2427]*kernel[7]+tmp[2428]*kernel[8];
				ans[2328]<=tmp[2227]*kernel[0]+tmp[2228]*kernel[1]+tmp[2229]*kernel[2]+tmp[2327]*kernel[3]+tmp[2328]*kernel[4]+tmp[2329]*kernel[5]+tmp[2427]*kernel[6]+tmp[2428]*kernel[7]+tmp[2429]*kernel[8];
				ans[2329]<=tmp[2228]*kernel[0]+tmp[2229]*kernel[1]+tmp[2230]*kernel[2]+tmp[2328]*kernel[3]+tmp[2329]*kernel[4]+tmp[2330]*kernel[5]+tmp[2428]*kernel[6]+tmp[2429]*kernel[7]+tmp[2430]*kernel[8];
				ans[2330]<=tmp[2229]*kernel[0]+tmp[2230]*kernel[1]+tmp[2231]*kernel[2]+tmp[2329]*kernel[3]+tmp[2330]*kernel[4]+tmp[2331]*kernel[5]+tmp[2429]*kernel[6]+tmp[2430]*kernel[7]+tmp[2431]*kernel[8];
				ans[2331]<=tmp[2230]*kernel[0]+tmp[2231]*kernel[1]+tmp[2232]*kernel[2]+tmp[2330]*kernel[3]+tmp[2331]*kernel[4]+tmp[2332]*kernel[5]+tmp[2430]*kernel[6]+tmp[2431]*kernel[7]+tmp[2432]*kernel[8];
				ans[2332]<=tmp[2231]*kernel[0]+tmp[2232]*kernel[1]+tmp[2233]*kernel[2]+tmp[2331]*kernel[3]+tmp[2332]*kernel[4]+tmp[2333]*kernel[5]+tmp[2431]*kernel[6]+tmp[2432]*kernel[7]+tmp[2433]*kernel[8];
				ans[2333]<=tmp[2232]*kernel[0]+tmp[2233]*kernel[1]+tmp[2234]*kernel[2]+tmp[2332]*kernel[3]+tmp[2333]*kernel[4]+tmp[2334]*kernel[5]+tmp[2432]*kernel[6]+tmp[2433]*kernel[7]+tmp[2434]*kernel[8];
				ans[2334]<=tmp[2233]*kernel[0]+tmp[2234]*kernel[1]+tmp[2235]*kernel[2]+tmp[2333]*kernel[3]+tmp[2334]*kernel[4]+tmp[2335]*kernel[5]+tmp[2433]*kernel[6]+tmp[2434]*kernel[7]+tmp[2435]*kernel[8];
				ans[2335]<=tmp[2234]*kernel[0]+tmp[2235]*kernel[1]+tmp[2236]*kernel[2]+tmp[2334]*kernel[3]+tmp[2335]*kernel[4]+tmp[2336]*kernel[5]+tmp[2434]*kernel[6]+tmp[2435]*kernel[7]+tmp[2436]*kernel[8];
				ans[2336]<=tmp[2235]*kernel[0]+tmp[2236]*kernel[1]+tmp[2237]*kernel[2]+tmp[2335]*kernel[3]+tmp[2336]*kernel[4]+tmp[2337]*kernel[5]+tmp[2435]*kernel[6]+tmp[2436]*kernel[7]+tmp[2437]*kernel[8];
				ans[2337]<=tmp[2236]*kernel[0]+tmp[2237]*kernel[1]+tmp[2238]*kernel[2]+tmp[2336]*kernel[3]+tmp[2337]*kernel[4]+tmp[2338]*kernel[5]+tmp[2436]*kernel[6]+tmp[2437]*kernel[7]+tmp[2438]*kernel[8];
				ans[2338]<=tmp[2237]*kernel[0]+tmp[2238]*kernel[1]+tmp[2239]*kernel[2]+tmp[2337]*kernel[3]+tmp[2338]*kernel[4]+tmp[2339]*kernel[5]+tmp[2437]*kernel[6]+tmp[2438]*kernel[7]+tmp[2439]*kernel[8];
				ans[2339]<=tmp[2238]*kernel[0]+tmp[2239]*kernel[1]+tmp[2240]*kernel[2]+tmp[2338]*kernel[3]+tmp[2339]*kernel[4]+tmp[2340]*kernel[5]+tmp[2438]*kernel[6]+tmp[2439]*kernel[7]+tmp[2440]*kernel[8];
				ans[2340]<=tmp[2239]*kernel[0]+tmp[2240]*kernel[1]+tmp[2241]*kernel[2]+tmp[2339]*kernel[3]+tmp[2340]*kernel[4]+tmp[2341]*kernel[5]+tmp[2439]*kernel[6]+tmp[2440]*kernel[7]+tmp[2441]*kernel[8];
				ans[2341]<=tmp[2240]*kernel[0]+tmp[2241]*kernel[1]+tmp[2242]*kernel[2]+tmp[2340]*kernel[3]+tmp[2341]*kernel[4]+tmp[2342]*kernel[5]+tmp[2440]*kernel[6]+tmp[2441]*kernel[7]+tmp[2442]*kernel[8];
				ans[2342]<=tmp[2241]*kernel[0]+tmp[2242]*kernel[1]+tmp[2243]*kernel[2]+tmp[2341]*kernel[3]+tmp[2342]*kernel[4]+tmp[2343]*kernel[5]+tmp[2441]*kernel[6]+tmp[2442]*kernel[7]+tmp[2443]*kernel[8];
				ans[2343]<=tmp[2242]*kernel[0]+tmp[2243]*kernel[1]+tmp[2244]*kernel[2]+tmp[2342]*kernel[3]+tmp[2343]*kernel[4]+tmp[2344]*kernel[5]+tmp[2442]*kernel[6]+tmp[2443]*kernel[7]+tmp[2444]*kernel[8];
				ans[2344]<=tmp[2243]*kernel[0]+tmp[2244]*kernel[1]+tmp[2245]*kernel[2]+tmp[2343]*kernel[3]+tmp[2344]*kernel[4]+tmp[2345]*kernel[5]+tmp[2443]*kernel[6]+tmp[2444]*kernel[7]+tmp[2445]*kernel[8];
				ans[2345]<=tmp[2244]*kernel[0]+tmp[2245]*kernel[1]+tmp[2246]*kernel[2]+tmp[2344]*kernel[3]+tmp[2345]*kernel[4]+tmp[2346]*kernel[5]+tmp[2444]*kernel[6]+tmp[2445]*kernel[7]+tmp[2446]*kernel[8];
				ans[2346]<=tmp[2245]*kernel[0]+tmp[2246]*kernel[1]+tmp[2247]*kernel[2]+tmp[2345]*kernel[3]+tmp[2346]*kernel[4]+tmp[2347]*kernel[5]+tmp[2445]*kernel[6]+tmp[2446]*kernel[7]+tmp[2447]*kernel[8];
				ans[2347]<=tmp[2246]*kernel[0]+tmp[2247]*kernel[1]+tmp[2248]*kernel[2]+tmp[2346]*kernel[3]+tmp[2347]*kernel[4]+tmp[2348]*kernel[5]+tmp[2446]*kernel[6]+tmp[2447]*kernel[7]+tmp[2448]*kernel[8];
				ans[2348]<=tmp[2247]*kernel[0]+tmp[2248]*kernel[1]+tmp[2249]*kernel[2]+tmp[2347]*kernel[3]+tmp[2348]*kernel[4]+tmp[2349]*kernel[5]+tmp[2447]*kernel[6]+tmp[2448]*kernel[7]+tmp[2449]*kernel[8];
				ans[2349]<=tmp[2248]*kernel[0]+tmp[2249]*kernel[1]+tmp[2250]*kernel[2]+tmp[2348]*kernel[3]+tmp[2349]*kernel[4]+tmp[2350]*kernel[5]+tmp[2448]*kernel[6]+tmp[2449]*kernel[7]+tmp[2450]*kernel[8];
				ans[2350]<=tmp[2249]*kernel[0]+tmp[2250]*kernel[1]+tmp[2251]*kernel[2]+tmp[2349]*kernel[3]+tmp[2350]*kernel[4]+tmp[2351]*kernel[5]+tmp[2449]*kernel[6]+tmp[2450]*kernel[7]+tmp[2451]*kernel[8];
				ans[2351]<=tmp[2250]*kernel[0]+tmp[2251]*kernel[1]+tmp[2252]*kernel[2]+tmp[2350]*kernel[3]+tmp[2351]*kernel[4]+tmp[2352]*kernel[5]+tmp[2450]*kernel[6]+tmp[2451]*kernel[7]+tmp[2452]*kernel[8];
				ans[2352]<=tmp[2251]*kernel[0]+tmp[2252]*kernel[1]+tmp[2253]*kernel[2]+tmp[2351]*kernel[3]+tmp[2352]*kernel[4]+tmp[2353]*kernel[5]+tmp[2451]*kernel[6]+tmp[2452]*kernel[7]+tmp[2453]*kernel[8];
				ans[2353]<=tmp[2252]*kernel[0]+tmp[2253]*kernel[1]+tmp[2254]*kernel[2]+tmp[2352]*kernel[3]+tmp[2353]*kernel[4]+tmp[2354]*kernel[5]+tmp[2452]*kernel[6]+tmp[2453]*kernel[7]+tmp[2454]*kernel[8];
				ans[2354]<=tmp[2253]*kernel[0]+tmp[2254]*kernel[1]+tmp[2255]*kernel[2]+tmp[2353]*kernel[3]+tmp[2354]*kernel[4]+tmp[2355]*kernel[5]+tmp[2453]*kernel[6]+tmp[2454]*kernel[7]+tmp[2455]*kernel[8];
				ans[2355]<=tmp[2254]*kernel[0]+tmp[2255]*kernel[1]+tmp[2256]*kernel[2]+tmp[2354]*kernel[3]+tmp[2355]*kernel[4]+tmp[2356]*kernel[5]+tmp[2454]*kernel[6]+tmp[2455]*kernel[7]+tmp[2456]*kernel[8];
				ans[2356]<=tmp[2255]*kernel[0]+tmp[2256]*kernel[1]+tmp[2257]*kernel[2]+tmp[2355]*kernel[3]+tmp[2356]*kernel[4]+tmp[2357]*kernel[5]+tmp[2455]*kernel[6]+tmp[2456]*kernel[7]+tmp[2457]*kernel[8];
				ans[2357]<=tmp[2256]*kernel[0]+tmp[2257]*kernel[1]+tmp[2258]*kernel[2]+tmp[2356]*kernel[3]+tmp[2357]*kernel[4]+tmp[2358]*kernel[5]+tmp[2456]*kernel[6]+tmp[2457]*kernel[7]+tmp[2458]*kernel[8];
				ans[2358]<=tmp[2257]*kernel[0]+tmp[2258]*kernel[1]+tmp[2259]*kernel[2]+tmp[2357]*kernel[3]+tmp[2358]*kernel[4]+tmp[2359]*kernel[5]+tmp[2457]*kernel[6]+tmp[2458]*kernel[7]+tmp[2459]*kernel[8];
				ans[2359]<=tmp[2258]*kernel[0]+tmp[2259]*kernel[1]+tmp[2260]*kernel[2]+tmp[2358]*kernel[3]+tmp[2359]*kernel[4]+tmp[2360]*kernel[5]+tmp[2458]*kernel[6]+tmp[2459]*kernel[7]+tmp[2460]*kernel[8];
				ans[2360]<=tmp[2259]*kernel[0]+tmp[2260]*kernel[1]+tmp[2261]*kernel[2]+tmp[2359]*kernel[3]+tmp[2360]*kernel[4]+tmp[2361]*kernel[5]+tmp[2459]*kernel[6]+tmp[2460]*kernel[7]+tmp[2461]*kernel[8];
				ans[2361]<=tmp[2260]*kernel[0]+tmp[2261]*kernel[1]+tmp[2262]*kernel[2]+tmp[2360]*kernel[3]+tmp[2361]*kernel[4]+tmp[2362]*kernel[5]+tmp[2460]*kernel[6]+tmp[2461]*kernel[7]+tmp[2462]*kernel[8];
				ans[2362]<=tmp[2261]*kernel[0]+tmp[2262]*kernel[1]+tmp[2263]*kernel[2]+tmp[2361]*kernel[3]+tmp[2362]*kernel[4]+tmp[2363]*kernel[5]+tmp[2461]*kernel[6]+tmp[2462]*kernel[7]+tmp[2463]*kernel[8];
				ans[2363]<=tmp[2262]*kernel[0]+tmp[2263]*kernel[1]+tmp[2264]*kernel[2]+tmp[2362]*kernel[3]+tmp[2363]*kernel[4]+tmp[2364]*kernel[5]+tmp[2462]*kernel[6]+tmp[2463]*kernel[7]+tmp[2464]*kernel[8];
				ans[2364]<=tmp[2263]*kernel[0]+tmp[2264]*kernel[1]+tmp[2265]*kernel[2]+tmp[2363]*kernel[3]+tmp[2364]*kernel[4]+tmp[2365]*kernel[5]+tmp[2463]*kernel[6]+tmp[2464]*kernel[7]+tmp[2465]*kernel[8];
				ans[2365]<=tmp[2264]*kernel[0]+tmp[2265]*kernel[1]+tmp[2266]*kernel[2]+tmp[2364]*kernel[3]+tmp[2365]*kernel[4]+tmp[2366]*kernel[5]+tmp[2464]*kernel[6]+tmp[2465]*kernel[7]+tmp[2466]*kernel[8];
				ans[2366]<=tmp[2265]*kernel[0]+tmp[2266]*kernel[1]+tmp[2267]*kernel[2]+tmp[2365]*kernel[3]+tmp[2366]*kernel[4]+tmp[2367]*kernel[5]+tmp[2465]*kernel[6]+tmp[2466]*kernel[7]+tmp[2467]*kernel[8];
				ans[2367]<=tmp[2266]*kernel[0]+tmp[2267]*kernel[1]+tmp[2268]*kernel[2]+tmp[2366]*kernel[3]+tmp[2367]*kernel[4]+tmp[2368]*kernel[5]+tmp[2466]*kernel[6]+tmp[2467]*kernel[7]+tmp[2468]*kernel[8];
				ans[2368]<=tmp[2267]*kernel[0]+tmp[2268]*kernel[1]+tmp[2269]*kernel[2]+tmp[2367]*kernel[3]+tmp[2368]*kernel[4]+tmp[2369]*kernel[5]+tmp[2467]*kernel[6]+tmp[2468]*kernel[7]+tmp[2469]*kernel[8];
				ans[2369]<=tmp[2268]*kernel[0]+tmp[2269]*kernel[1]+tmp[2270]*kernel[2]+tmp[2368]*kernel[3]+tmp[2369]*kernel[4]+tmp[2370]*kernel[5]+tmp[2468]*kernel[6]+tmp[2469]*kernel[7]+tmp[2470]*kernel[8];
				ans[2370]<=tmp[2269]*kernel[0]+tmp[2270]*kernel[1]+tmp[2271]*kernel[2]+tmp[2369]*kernel[3]+tmp[2370]*kernel[4]+tmp[2371]*kernel[5]+tmp[2469]*kernel[6]+tmp[2470]*kernel[7]+tmp[2471]*kernel[8];
				ans[2371]<=tmp[2270]*kernel[0]+tmp[2271]*kernel[1]+tmp[2272]*kernel[2]+tmp[2370]*kernel[3]+tmp[2371]*kernel[4]+tmp[2372]*kernel[5]+tmp[2470]*kernel[6]+tmp[2471]*kernel[7]+tmp[2472]*kernel[8];
				ans[2372]<=tmp[2271]*kernel[0]+tmp[2272]*kernel[1]+tmp[2273]*kernel[2]+tmp[2371]*kernel[3]+tmp[2372]*kernel[4]+tmp[2373]*kernel[5]+tmp[2471]*kernel[6]+tmp[2472]*kernel[7]+tmp[2473]*kernel[8];
				ans[2373]<=tmp[2272]*kernel[0]+tmp[2273]*kernel[1]+tmp[2274]*kernel[2]+tmp[2372]*kernel[3]+tmp[2373]*kernel[4]+tmp[2374]*kernel[5]+tmp[2472]*kernel[6]+tmp[2473]*kernel[7]+tmp[2474]*kernel[8];
				ans[2374]<=tmp[2273]*kernel[0]+tmp[2274]*kernel[1]+tmp[2275]*kernel[2]+tmp[2373]*kernel[3]+tmp[2374]*kernel[4]+tmp[2375]*kernel[5]+tmp[2473]*kernel[6]+tmp[2474]*kernel[7]+tmp[2475]*kernel[8];
				ans[2375]<=tmp[2274]*kernel[0]+tmp[2275]*kernel[1]+tmp[2276]*kernel[2]+tmp[2374]*kernel[3]+tmp[2375]*kernel[4]+tmp[2376]*kernel[5]+tmp[2474]*kernel[6]+tmp[2475]*kernel[7]+tmp[2476]*kernel[8];
				ans[2376]<=tmp[2275]*kernel[0]+tmp[2276]*kernel[1]+tmp[2277]*kernel[2]+tmp[2375]*kernel[3]+tmp[2376]*kernel[4]+tmp[2377]*kernel[5]+tmp[2475]*kernel[6]+tmp[2476]*kernel[7]+tmp[2477]*kernel[8];
				ans[2377]<=tmp[2276]*kernel[0]+tmp[2277]*kernel[1]+tmp[2278]*kernel[2]+tmp[2376]*kernel[3]+tmp[2377]*kernel[4]+tmp[2378]*kernel[5]+tmp[2476]*kernel[6]+tmp[2477]*kernel[7]+tmp[2478]*kernel[8];
				ans[2378]<=tmp[2277]*kernel[0]+tmp[2278]*kernel[1]+tmp[2279]*kernel[2]+tmp[2377]*kernel[3]+tmp[2378]*kernel[4]+tmp[2379]*kernel[5]+tmp[2477]*kernel[6]+tmp[2478]*kernel[7]+tmp[2479]*kernel[8];
				ans[2379]<=tmp[2278]*kernel[0]+tmp[2279]*kernel[1]+tmp[2280]*kernel[2]+tmp[2378]*kernel[3]+tmp[2379]*kernel[4]+tmp[2380]*kernel[5]+tmp[2478]*kernel[6]+tmp[2479]*kernel[7]+tmp[2480]*kernel[8];
				ans[2380]<=tmp[2279]*kernel[0]+tmp[2280]*kernel[1]+tmp[2281]*kernel[2]+tmp[2379]*kernel[3]+tmp[2380]*kernel[4]+tmp[2381]*kernel[5]+tmp[2479]*kernel[6]+tmp[2480]*kernel[7]+tmp[2481]*kernel[8];
				ans[2381]<=tmp[2280]*kernel[0]+tmp[2281]*kernel[1]+tmp[2282]*kernel[2]+tmp[2380]*kernel[3]+tmp[2381]*kernel[4]+tmp[2382]*kernel[5]+tmp[2480]*kernel[6]+tmp[2481]*kernel[7]+tmp[2482]*kernel[8];
				ans[2382]<=tmp[2281]*kernel[0]+tmp[2282]*kernel[1]+tmp[2283]*kernel[2]+tmp[2381]*kernel[3]+tmp[2382]*kernel[4]+tmp[2383]*kernel[5]+tmp[2481]*kernel[6]+tmp[2482]*kernel[7]+tmp[2483]*kernel[8];
				ans[2383]<=tmp[2282]*kernel[0]+tmp[2283]*kernel[1]+tmp[2284]*kernel[2]+tmp[2382]*kernel[3]+tmp[2383]*kernel[4]+tmp[2384]*kernel[5]+tmp[2482]*kernel[6]+tmp[2483]*kernel[7]+tmp[2484]*kernel[8];
				ans[2384]<=tmp[2283]*kernel[0]+tmp[2284]*kernel[1]+tmp[2285]*kernel[2]+tmp[2383]*kernel[3]+tmp[2384]*kernel[4]+tmp[2385]*kernel[5]+tmp[2483]*kernel[6]+tmp[2484]*kernel[7]+tmp[2485]*kernel[8];
				ans[2385]<=tmp[2284]*kernel[0]+tmp[2285]*kernel[1]+tmp[2286]*kernel[2]+tmp[2384]*kernel[3]+tmp[2385]*kernel[4]+tmp[2386]*kernel[5]+tmp[2484]*kernel[6]+tmp[2485]*kernel[7]+tmp[2486]*kernel[8];
				ans[2386]<=tmp[2285]*kernel[0]+tmp[2286]*kernel[1]+tmp[2287]*kernel[2]+tmp[2385]*kernel[3]+tmp[2386]*kernel[4]+tmp[2387]*kernel[5]+tmp[2485]*kernel[6]+tmp[2486]*kernel[7]+tmp[2487]*kernel[8];
				ans[2387]<=tmp[2286]*kernel[0]+tmp[2287]*kernel[1]+tmp[2288]*kernel[2]+tmp[2386]*kernel[3]+tmp[2387]*kernel[4]+tmp[2388]*kernel[5]+tmp[2486]*kernel[6]+tmp[2487]*kernel[7]+tmp[2488]*kernel[8];
				ans[2388]<=tmp[2287]*kernel[0]+tmp[2288]*kernel[1]+tmp[2289]*kernel[2]+tmp[2387]*kernel[3]+tmp[2388]*kernel[4]+tmp[2389]*kernel[5]+tmp[2487]*kernel[6]+tmp[2488]*kernel[7]+tmp[2489]*kernel[8];
				ans[2389]<=tmp[2288]*kernel[0]+tmp[2289]*kernel[1]+tmp[2290]*kernel[2]+tmp[2388]*kernel[3]+tmp[2389]*kernel[4]+tmp[2390]*kernel[5]+tmp[2488]*kernel[6]+tmp[2489]*kernel[7]+tmp[2490]*kernel[8];
				ans[2390]<=tmp[2289]*kernel[0]+tmp[2290]*kernel[1]+tmp[2291]*kernel[2]+tmp[2389]*kernel[3]+tmp[2390]*kernel[4]+tmp[2391]*kernel[5]+tmp[2489]*kernel[6]+tmp[2490]*kernel[7]+tmp[2491]*kernel[8];
				ans[2391]<=tmp[2290]*kernel[0]+tmp[2291]*kernel[1]+tmp[2292]*kernel[2]+tmp[2390]*kernel[3]+tmp[2391]*kernel[4]+tmp[2392]*kernel[5]+tmp[2490]*kernel[6]+tmp[2491]*kernel[7]+tmp[2492]*kernel[8];
				ans[2392]<=tmp[2291]*kernel[0]+tmp[2292]*kernel[1]+tmp[2293]*kernel[2]+tmp[2391]*kernel[3]+tmp[2392]*kernel[4]+tmp[2393]*kernel[5]+tmp[2491]*kernel[6]+tmp[2492]*kernel[7]+tmp[2493]*kernel[8];
				ans[2393]<=tmp[2292]*kernel[0]+tmp[2293]*kernel[1]+tmp[2294]*kernel[2]+tmp[2392]*kernel[3]+tmp[2393]*kernel[4]+tmp[2394]*kernel[5]+tmp[2492]*kernel[6]+tmp[2493]*kernel[7]+tmp[2494]*kernel[8];
				ans[2394]<=tmp[2293]*kernel[0]+tmp[2294]*kernel[1]+tmp[2295]*kernel[2]+tmp[2393]*kernel[3]+tmp[2394]*kernel[4]+tmp[2395]*kernel[5]+tmp[2493]*kernel[6]+tmp[2494]*kernel[7]+tmp[2495]*kernel[8];
				ans[2395]<=tmp[2294]*kernel[0]+tmp[2295]*kernel[1]+tmp[2296]*kernel[2]+tmp[2394]*kernel[3]+tmp[2395]*kernel[4]+tmp[2396]*kernel[5]+tmp[2494]*kernel[6]+tmp[2495]*kernel[7]+tmp[2496]*kernel[8];
				ans[2396]<=tmp[2295]*kernel[0]+tmp[2296]*kernel[1]+tmp[2297]*kernel[2]+tmp[2395]*kernel[3]+tmp[2396]*kernel[4]+tmp[2397]*kernel[5]+tmp[2495]*kernel[6]+tmp[2496]*kernel[7]+tmp[2497]*kernel[8];
				ans[2397]<=tmp[2296]*kernel[0]+tmp[2297]*kernel[1]+tmp[2298]*kernel[2]+tmp[2396]*kernel[3]+tmp[2397]*kernel[4]+tmp[2398]*kernel[5]+tmp[2496]*kernel[6]+tmp[2497]*kernel[7]+tmp[2498]*kernel[8];
				ans[2398]<=tmp[2297]*kernel[0]+tmp[2298]*kernel[1]+tmp[2299]*kernel[2]+tmp[2397]*kernel[3]+tmp[2398]*kernel[4]+tmp[2399]*kernel[5]+tmp[2497]*kernel[6]+tmp[2498]*kernel[7]+tmp[2499]*kernel[8];
				ans[2399]<=tmp[2298]*kernel[0]+tmp[2299]*kernel[1]+tmp[2398]*kernel[3]+tmp[2399]*kernel[4]+tmp[2498]*kernel[6]+tmp[2499]*kernel[7];
				ans[2400]<=tmp[2300]*kernel[1]+tmp[2301]*kernel[2]+tmp[2400]*kernel[4]+tmp[2401]*kernel[5]+tmp[2500]*kernel[7]+tmp[2501]*kernel[8];
				ans[2401]<=tmp[2300]*kernel[0]+tmp[2301]*kernel[1]+tmp[2302]*kernel[2]+tmp[2400]*kernel[3]+tmp[2401]*kernel[4]+tmp[2402]*kernel[5]+tmp[2500]*kernel[6]+tmp[2501]*kernel[7]+tmp[2502]*kernel[8];
				ans[2402]<=tmp[2301]*kernel[0]+tmp[2302]*kernel[1]+tmp[2303]*kernel[2]+tmp[2401]*kernel[3]+tmp[2402]*kernel[4]+tmp[2403]*kernel[5]+tmp[2501]*kernel[6]+tmp[2502]*kernel[7]+tmp[2503]*kernel[8];
				ans[2403]<=tmp[2302]*kernel[0]+tmp[2303]*kernel[1]+tmp[2304]*kernel[2]+tmp[2402]*kernel[3]+tmp[2403]*kernel[4]+tmp[2404]*kernel[5]+tmp[2502]*kernel[6]+tmp[2503]*kernel[7]+tmp[2504]*kernel[8];
				ans[2404]<=tmp[2303]*kernel[0]+tmp[2304]*kernel[1]+tmp[2305]*kernel[2]+tmp[2403]*kernel[3]+tmp[2404]*kernel[4]+tmp[2405]*kernel[5]+tmp[2503]*kernel[6]+tmp[2504]*kernel[7]+tmp[2505]*kernel[8];
				ans[2405]<=tmp[2304]*kernel[0]+tmp[2305]*kernel[1]+tmp[2306]*kernel[2]+tmp[2404]*kernel[3]+tmp[2405]*kernel[4]+tmp[2406]*kernel[5]+tmp[2504]*kernel[6]+tmp[2505]*kernel[7]+tmp[2506]*kernel[8];
				ans[2406]<=tmp[2305]*kernel[0]+tmp[2306]*kernel[1]+tmp[2307]*kernel[2]+tmp[2405]*kernel[3]+tmp[2406]*kernel[4]+tmp[2407]*kernel[5]+tmp[2505]*kernel[6]+tmp[2506]*kernel[7]+tmp[2507]*kernel[8];
				ans[2407]<=tmp[2306]*kernel[0]+tmp[2307]*kernel[1]+tmp[2308]*kernel[2]+tmp[2406]*kernel[3]+tmp[2407]*kernel[4]+tmp[2408]*kernel[5]+tmp[2506]*kernel[6]+tmp[2507]*kernel[7]+tmp[2508]*kernel[8];
				ans[2408]<=tmp[2307]*kernel[0]+tmp[2308]*kernel[1]+tmp[2309]*kernel[2]+tmp[2407]*kernel[3]+tmp[2408]*kernel[4]+tmp[2409]*kernel[5]+tmp[2507]*kernel[6]+tmp[2508]*kernel[7]+tmp[2509]*kernel[8];
				ans[2409]<=tmp[2308]*kernel[0]+tmp[2309]*kernel[1]+tmp[2310]*kernel[2]+tmp[2408]*kernel[3]+tmp[2409]*kernel[4]+tmp[2410]*kernel[5]+tmp[2508]*kernel[6]+tmp[2509]*kernel[7]+tmp[2510]*kernel[8];
				ans[2410]<=tmp[2309]*kernel[0]+tmp[2310]*kernel[1]+tmp[2311]*kernel[2]+tmp[2409]*kernel[3]+tmp[2410]*kernel[4]+tmp[2411]*kernel[5]+tmp[2509]*kernel[6]+tmp[2510]*kernel[7]+tmp[2511]*kernel[8];
				ans[2411]<=tmp[2310]*kernel[0]+tmp[2311]*kernel[1]+tmp[2312]*kernel[2]+tmp[2410]*kernel[3]+tmp[2411]*kernel[4]+tmp[2412]*kernel[5]+tmp[2510]*kernel[6]+tmp[2511]*kernel[7]+tmp[2512]*kernel[8];
				ans[2412]<=tmp[2311]*kernel[0]+tmp[2312]*kernel[1]+tmp[2313]*kernel[2]+tmp[2411]*kernel[3]+tmp[2412]*kernel[4]+tmp[2413]*kernel[5]+tmp[2511]*kernel[6]+tmp[2512]*kernel[7]+tmp[2513]*kernel[8];
				ans[2413]<=tmp[2312]*kernel[0]+tmp[2313]*kernel[1]+tmp[2314]*kernel[2]+tmp[2412]*kernel[3]+tmp[2413]*kernel[4]+tmp[2414]*kernel[5]+tmp[2512]*kernel[6]+tmp[2513]*kernel[7]+tmp[2514]*kernel[8];
				ans[2414]<=tmp[2313]*kernel[0]+tmp[2314]*kernel[1]+tmp[2315]*kernel[2]+tmp[2413]*kernel[3]+tmp[2414]*kernel[4]+tmp[2415]*kernel[5]+tmp[2513]*kernel[6]+tmp[2514]*kernel[7]+tmp[2515]*kernel[8];
				ans[2415]<=tmp[2314]*kernel[0]+tmp[2315]*kernel[1]+tmp[2316]*kernel[2]+tmp[2414]*kernel[3]+tmp[2415]*kernel[4]+tmp[2416]*kernel[5]+tmp[2514]*kernel[6]+tmp[2515]*kernel[7]+tmp[2516]*kernel[8];
				ans[2416]<=tmp[2315]*kernel[0]+tmp[2316]*kernel[1]+tmp[2317]*kernel[2]+tmp[2415]*kernel[3]+tmp[2416]*kernel[4]+tmp[2417]*kernel[5]+tmp[2515]*kernel[6]+tmp[2516]*kernel[7]+tmp[2517]*kernel[8];
				ans[2417]<=tmp[2316]*kernel[0]+tmp[2317]*kernel[1]+tmp[2318]*kernel[2]+tmp[2416]*kernel[3]+tmp[2417]*kernel[4]+tmp[2418]*kernel[5]+tmp[2516]*kernel[6]+tmp[2517]*kernel[7]+tmp[2518]*kernel[8];
				ans[2418]<=tmp[2317]*kernel[0]+tmp[2318]*kernel[1]+tmp[2319]*kernel[2]+tmp[2417]*kernel[3]+tmp[2418]*kernel[4]+tmp[2419]*kernel[5]+tmp[2517]*kernel[6]+tmp[2518]*kernel[7]+tmp[2519]*kernel[8];
				ans[2419]<=tmp[2318]*kernel[0]+tmp[2319]*kernel[1]+tmp[2320]*kernel[2]+tmp[2418]*kernel[3]+tmp[2419]*kernel[4]+tmp[2420]*kernel[5]+tmp[2518]*kernel[6]+tmp[2519]*kernel[7]+tmp[2520]*kernel[8];
				ans[2420]<=tmp[2319]*kernel[0]+tmp[2320]*kernel[1]+tmp[2321]*kernel[2]+tmp[2419]*kernel[3]+tmp[2420]*kernel[4]+tmp[2421]*kernel[5]+tmp[2519]*kernel[6]+tmp[2520]*kernel[7]+tmp[2521]*kernel[8];
				ans[2421]<=tmp[2320]*kernel[0]+tmp[2321]*kernel[1]+tmp[2322]*kernel[2]+tmp[2420]*kernel[3]+tmp[2421]*kernel[4]+tmp[2422]*kernel[5]+tmp[2520]*kernel[6]+tmp[2521]*kernel[7]+tmp[2522]*kernel[8];
				ans[2422]<=tmp[2321]*kernel[0]+tmp[2322]*kernel[1]+tmp[2323]*kernel[2]+tmp[2421]*kernel[3]+tmp[2422]*kernel[4]+tmp[2423]*kernel[5]+tmp[2521]*kernel[6]+tmp[2522]*kernel[7]+tmp[2523]*kernel[8];
				ans[2423]<=tmp[2322]*kernel[0]+tmp[2323]*kernel[1]+tmp[2324]*kernel[2]+tmp[2422]*kernel[3]+tmp[2423]*kernel[4]+tmp[2424]*kernel[5]+tmp[2522]*kernel[6]+tmp[2523]*kernel[7]+tmp[2524]*kernel[8];
				ans[2424]<=tmp[2323]*kernel[0]+tmp[2324]*kernel[1]+tmp[2325]*kernel[2]+tmp[2423]*kernel[3]+tmp[2424]*kernel[4]+tmp[2425]*kernel[5]+tmp[2523]*kernel[6]+tmp[2524]*kernel[7]+tmp[2525]*kernel[8];
				ans[2425]<=tmp[2324]*kernel[0]+tmp[2325]*kernel[1]+tmp[2326]*kernel[2]+tmp[2424]*kernel[3]+tmp[2425]*kernel[4]+tmp[2426]*kernel[5]+tmp[2524]*kernel[6]+tmp[2525]*kernel[7]+tmp[2526]*kernel[8];
				ans[2426]<=tmp[2325]*kernel[0]+tmp[2326]*kernel[1]+tmp[2327]*kernel[2]+tmp[2425]*kernel[3]+tmp[2426]*kernel[4]+tmp[2427]*kernel[5]+tmp[2525]*kernel[6]+tmp[2526]*kernel[7]+tmp[2527]*kernel[8];
				ans[2427]<=tmp[2326]*kernel[0]+tmp[2327]*kernel[1]+tmp[2328]*kernel[2]+tmp[2426]*kernel[3]+tmp[2427]*kernel[4]+tmp[2428]*kernel[5]+tmp[2526]*kernel[6]+tmp[2527]*kernel[7]+tmp[2528]*kernel[8];
				ans[2428]<=tmp[2327]*kernel[0]+tmp[2328]*kernel[1]+tmp[2329]*kernel[2]+tmp[2427]*kernel[3]+tmp[2428]*kernel[4]+tmp[2429]*kernel[5]+tmp[2527]*kernel[6]+tmp[2528]*kernel[7]+tmp[2529]*kernel[8];
				ans[2429]<=tmp[2328]*kernel[0]+tmp[2329]*kernel[1]+tmp[2330]*kernel[2]+tmp[2428]*kernel[3]+tmp[2429]*kernel[4]+tmp[2430]*kernel[5]+tmp[2528]*kernel[6]+tmp[2529]*kernel[7]+tmp[2530]*kernel[8];
				ans[2430]<=tmp[2329]*kernel[0]+tmp[2330]*kernel[1]+tmp[2331]*kernel[2]+tmp[2429]*kernel[3]+tmp[2430]*kernel[4]+tmp[2431]*kernel[5]+tmp[2529]*kernel[6]+tmp[2530]*kernel[7]+tmp[2531]*kernel[8];
				ans[2431]<=tmp[2330]*kernel[0]+tmp[2331]*kernel[1]+tmp[2332]*kernel[2]+tmp[2430]*kernel[3]+tmp[2431]*kernel[4]+tmp[2432]*kernel[5]+tmp[2530]*kernel[6]+tmp[2531]*kernel[7]+tmp[2532]*kernel[8];
				ans[2432]<=tmp[2331]*kernel[0]+tmp[2332]*kernel[1]+tmp[2333]*kernel[2]+tmp[2431]*kernel[3]+tmp[2432]*kernel[4]+tmp[2433]*kernel[5]+tmp[2531]*kernel[6]+tmp[2532]*kernel[7]+tmp[2533]*kernel[8];
				ans[2433]<=tmp[2332]*kernel[0]+tmp[2333]*kernel[1]+tmp[2334]*kernel[2]+tmp[2432]*kernel[3]+tmp[2433]*kernel[4]+tmp[2434]*kernel[5]+tmp[2532]*kernel[6]+tmp[2533]*kernel[7]+tmp[2534]*kernel[8];
				ans[2434]<=tmp[2333]*kernel[0]+tmp[2334]*kernel[1]+tmp[2335]*kernel[2]+tmp[2433]*kernel[3]+tmp[2434]*kernel[4]+tmp[2435]*kernel[5]+tmp[2533]*kernel[6]+tmp[2534]*kernel[7]+tmp[2535]*kernel[8];
				ans[2435]<=tmp[2334]*kernel[0]+tmp[2335]*kernel[1]+tmp[2336]*kernel[2]+tmp[2434]*kernel[3]+tmp[2435]*kernel[4]+tmp[2436]*kernel[5]+tmp[2534]*kernel[6]+tmp[2535]*kernel[7]+tmp[2536]*kernel[8];
				ans[2436]<=tmp[2335]*kernel[0]+tmp[2336]*kernel[1]+tmp[2337]*kernel[2]+tmp[2435]*kernel[3]+tmp[2436]*kernel[4]+tmp[2437]*kernel[5]+tmp[2535]*kernel[6]+tmp[2536]*kernel[7]+tmp[2537]*kernel[8];
				ans[2437]<=tmp[2336]*kernel[0]+tmp[2337]*kernel[1]+tmp[2338]*kernel[2]+tmp[2436]*kernel[3]+tmp[2437]*kernel[4]+tmp[2438]*kernel[5]+tmp[2536]*kernel[6]+tmp[2537]*kernel[7]+tmp[2538]*kernel[8];
				ans[2438]<=tmp[2337]*kernel[0]+tmp[2338]*kernel[1]+tmp[2339]*kernel[2]+tmp[2437]*kernel[3]+tmp[2438]*kernel[4]+tmp[2439]*kernel[5]+tmp[2537]*kernel[6]+tmp[2538]*kernel[7]+tmp[2539]*kernel[8];
				ans[2439]<=tmp[2338]*kernel[0]+tmp[2339]*kernel[1]+tmp[2340]*kernel[2]+tmp[2438]*kernel[3]+tmp[2439]*kernel[4]+tmp[2440]*kernel[5]+tmp[2538]*kernel[6]+tmp[2539]*kernel[7]+tmp[2540]*kernel[8];
				ans[2440]<=tmp[2339]*kernel[0]+tmp[2340]*kernel[1]+tmp[2341]*kernel[2]+tmp[2439]*kernel[3]+tmp[2440]*kernel[4]+tmp[2441]*kernel[5]+tmp[2539]*kernel[6]+tmp[2540]*kernel[7]+tmp[2541]*kernel[8];
				ans[2441]<=tmp[2340]*kernel[0]+tmp[2341]*kernel[1]+tmp[2342]*kernel[2]+tmp[2440]*kernel[3]+tmp[2441]*kernel[4]+tmp[2442]*kernel[5]+tmp[2540]*kernel[6]+tmp[2541]*kernel[7]+tmp[2542]*kernel[8];
				ans[2442]<=tmp[2341]*kernel[0]+tmp[2342]*kernel[1]+tmp[2343]*kernel[2]+tmp[2441]*kernel[3]+tmp[2442]*kernel[4]+tmp[2443]*kernel[5]+tmp[2541]*kernel[6]+tmp[2542]*kernel[7]+tmp[2543]*kernel[8];
				ans[2443]<=tmp[2342]*kernel[0]+tmp[2343]*kernel[1]+tmp[2344]*kernel[2]+tmp[2442]*kernel[3]+tmp[2443]*kernel[4]+tmp[2444]*kernel[5]+tmp[2542]*kernel[6]+tmp[2543]*kernel[7]+tmp[2544]*kernel[8];
				ans[2444]<=tmp[2343]*kernel[0]+tmp[2344]*kernel[1]+tmp[2345]*kernel[2]+tmp[2443]*kernel[3]+tmp[2444]*kernel[4]+tmp[2445]*kernel[5]+tmp[2543]*kernel[6]+tmp[2544]*kernel[7]+tmp[2545]*kernel[8];
				ans[2445]<=tmp[2344]*kernel[0]+tmp[2345]*kernel[1]+tmp[2346]*kernel[2]+tmp[2444]*kernel[3]+tmp[2445]*kernel[4]+tmp[2446]*kernel[5]+tmp[2544]*kernel[6]+tmp[2545]*kernel[7]+tmp[2546]*kernel[8];
				ans[2446]<=tmp[2345]*kernel[0]+tmp[2346]*kernel[1]+tmp[2347]*kernel[2]+tmp[2445]*kernel[3]+tmp[2446]*kernel[4]+tmp[2447]*kernel[5]+tmp[2545]*kernel[6]+tmp[2546]*kernel[7]+tmp[2547]*kernel[8];
				ans[2447]<=tmp[2346]*kernel[0]+tmp[2347]*kernel[1]+tmp[2348]*kernel[2]+tmp[2446]*kernel[3]+tmp[2447]*kernel[4]+tmp[2448]*kernel[5]+tmp[2546]*kernel[6]+tmp[2547]*kernel[7]+tmp[2548]*kernel[8];
				ans[2448]<=tmp[2347]*kernel[0]+tmp[2348]*kernel[1]+tmp[2349]*kernel[2]+tmp[2447]*kernel[3]+tmp[2448]*kernel[4]+tmp[2449]*kernel[5]+tmp[2547]*kernel[6]+tmp[2548]*kernel[7]+tmp[2549]*kernel[8];
				ans[2449]<=tmp[2348]*kernel[0]+tmp[2349]*kernel[1]+tmp[2350]*kernel[2]+tmp[2448]*kernel[3]+tmp[2449]*kernel[4]+tmp[2450]*kernel[5]+tmp[2548]*kernel[6]+tmp[2549]*kernel[7]+tmp[2550]*kernel[8];
				ans[2450]<=tmp[2349]*kernel[0]+tmp[2350]*kernel[1]+tmp[2351]*kernel[2]+tmp[2449]*kernel[3]+tmp[2450]*kernel[4]+tmp[2451]*kernel[5]+tmp[2549]*kernel[6]+tmp[2550]*kernel[7]+tmp[2551]*kernel[8];
				ans[2451]<=tmp[2350]*kernel[0]+tmp[2351]*kernel[1]+tmp[2352]*kernel[2]+tmp[2450]*kernel[3]+tmp[2451]*kernel[4]+tmp[2452]*kernel[5]+tmp[2550]*kernel[6]+tmp[2551]*kernel[7]+tmp[2552]*kernel[8];
				ans[2452]<=tmp[2351]*kernel[0]+tmp[2352]*kernel[1]+tmp[2353]*kernel[2]+tmp[2451]*kernel[3]+tmp[2452]*kernel[4]+tmp[2453]*kernel[5]+tmp[2551]*kernel[6]+tmp[2552]*kernel[7]+tmp[2553]*kernel[8];
				ans[2453]<=tmp[2352]*kernel[0]+tmp[2353]*kernel[1]+tmp[2354]*kernel[2]+tmp[2452]*kernel[3]+tmp[2453]*kernel[4]+tmp[2454]*kernel[5]+tmp[2552]*kernel[6]+tmp[2553]*kernel[7]+tmp[2554]*kernel[8];
				ans[2454]<=tmp[2353]*kernel[0]+tmp[2354]*kernel[1]+tmp[2355]*kernel[2]+tmp[2453]*kernel[3]+tmp[2454]*kernel[4]+tmp[2455]*kernel[5]+tmp[2553]*kernel[6]+tmp[2554]*kernel[7]+tmp[2555]*kernel[8];
				ans[2455]<=tmp[2354]*kernel[0]+tmp[2355]*kernel[1]+tmp[2356]*kernel[2]+tmp[2454]*kernel[3]+tmp[2455]*kernel[4]+tmp[2456]*kernel[5]+tmp[2554]*kernel[6]+tmp[2555]*kernel[7]+tmp[2556]*kernel[8];
				ans[2456]<=tmp[2355]*kernel[0]+tmp[2356]*kernel[1]+tmp[2357]*kernel[2]+tmp[2455]*kernel[3]+tmp[2456]*kernel[4]+tmp[2457]*kernel[5]+tmp[2555]*kernel[6]+tmp[2556]*kernel[7]+tmp[2557]*kernel[8];
				ans[2457]<=tmp[2356]*kernel[0]+tmp[2357]*kernel[1]+tmp[2358]*kernel[2]+tmp[2456]*kernel[3]+tmp[2457]*kernel[4]+tmp[2458]*kernel[5]+tmp[2556]*kernel[6]+tmp[2557]*kernel[7]+tmp[2558]*kernel[8];
				ans[2458]<=tmp[2357]*kernel[0]+tmp[2358]*kernel[1]+tmp[2359]*kernel[2]+tmp[2457]*kernel[3]+tmp[2458]*kernel[4]+tmp[2459]*kernel[5]+tmp[2557]*kernel[6]+tmp[2558]*kernel[7]+tmp[2559]*kernel[8];
				ans[2459]<=tmp[2358]*kernel[0]+tmp[2359]*kernel[1]+tmp[2360]*kernel[2]+tmp[2458]*kernel[3]+tmp[2459]*kernel[4]+tmp[2460]*kernel[5]+tmp[2558]*kernel[6]+tmp[2559]*kernel[7]+tmp[2560]*kernel[8];
				ans[2460]<=tmp[2359]*kernel[0]+tmp[2360]*kernel[1]+tmp[2361]*kernel[2]+tmp[2459]*kernel[3]+tmp[2460]*kernel[4]+tmp[2461]*kernel[5]+tmp[2559]*kernel[6]+tmp[2560]*kernel[7]+tmp[2561]*kernel[8];
				ans[2461]<=tmp[2360]*kernel[0]+tmp[2361]*kernel[1]+tmp[2362]*kernel[2]+tmp[2460]*kernel[3]+tmp[2461]*kernel[4]+tmp[2462]*kernel[5]+tmp[2560]*kernel[6]+tmp[2561]*kernel[7]+tmp[2562]*kernel[8];
				ans[2462]<=tmp[2361]*kernel[0]+tmp[2362]*kernel[1]+tmp[2363]*kernel[2]+tmp[2461]*kernel[3]+tmp[2462]*kernel[4]+tmp[2463]*kernel[5]+tmp[2561]*kernel[6]+tmp[2562]*kernel[7]+tmp[2563]*kernel[8];
				ans[2463]<=tmp[2362]*kernel[0]+tmp[2363]*kernel[1]+tmp[2364]*kernel[2]+tmp[2462]*kernel[3]+tmp[2463]*kernel[4]+tmp[2464]*kernel[5]+tmp[2562]*kernel[6]+tmp[2563]*kernel[7]+tmp[2564]*kernel[8];
				ans[2464]<=tmp[2363]*kernel[0]+tmp[2364]*kernel[1]+tmp[2365]*kernel[2]+tmp[2463]*kernel[3]+tmp[2464]*kernel[4]+tmp[2465]*kernel[5]+tmp[2563]*kernel[6]+tmp[2564]*kernel[7]+tmp[2565]*kernel[8];
				ans[2465]<=tmp[2364]*kernel[0]+tmp[2365]*kernel[1]+tmp[2366]*kernel[2]+tmp[2464]*kernel[3]+tmp[2465]*kernel[4]+tmp[2466]*kernel[5]+tmp[2564]*kernel[6]+tmp[2565]*kernel[7]+tmp[2566]*kernel[8];
				ans[2466]<=tmp[2365]*kernel[0]+tmp[2366]*kernel[1]+tmp[2367]*kernel[2]+tmp[2465]*kernel[3]+tmp[2466]*kernel[4]+tmp[2467]*kernel[5]+tmp[2565]*kernel[6]+tmp[2566]*kernel[7]+tmp[2567]*kernel[8];
				ans[2467]<=tmp[2366]*kernel[0]+tmp[2367]*kernel[1]+tmp[2368]*kernel[2]+tmp[2466]*kernel[3]+tmp[2467]*kernel[4]+tmp[2468]*kernel[5]+tmp[2566]*kernel[6]+tmp[2567]*kernel[7]+tmp[2568]*kernel[8];
				ans[2468]<=tmp[2367]*kernel[0]+tmp[2368]*kernel[1]+tmp[2369]*kernel[2]+tmp[2467]*kernel[3]+tmp[2468]*kernel[4]+tmp[2469]*kernel[5]+tmp[2567]*kernel[6]+tmp[2568]*kernel[7]+tmp[2569]*kernel[8];
				ans[2469]<=tmp[2368]*kernel[0]+tmp[2369]*kernel[1]+tmp[2370]*kernel[2]+tmp[2468]*kernel[3]+tmp[2469]*kernel[4]+tmp[2470]*kernel[5]+tmp[2568]*kernel[6]+tmp[2569]*kernel[7]+tmp[2570]*kernel[8];
				ans[2470]<=tmp[2369]*kernel[0]+tmp[2370]*kernel[1]+tmp[2371]*kernel[2]+tmp[2469]*kernel[3]+tmp[2470]*kernel[4]+tmp[2471]*kernel[5]+tmp[2569]*kernel[6]+tmp[2570]*kernel[7]+tmp[2571]*kernel[8];
				ans[2471]<=tmp[2370]*kernel[0]+tmp[2371]*kernel[1]+tmp[2372]*kernel[2]+tmp[2470]*kernel[3]+tmp[2471]*kernel[4]+tmp[2472]*kernel[5]+tmp[2570]*kernel[6]+tmp[2571]*kernel[7]+tmp[2572]*kernel[8];
				ans[2472]<=tmp[2371]*kernel[0]+tmp[2372]*kernel[1]+tmp[2373]*kernel[2]+tmp[2471]*kernel[3]+tmp[2472]*kernel[4]+tmp[2473]*kernel[5]+tmp[2571]*kernel[6]+tmp[2572]*kernel[7]+tmp[2573]*kernel[8];
				ans[2473]<=tmp[2372]*kernel[0]+tmp[2373]*kernel[1]+tmp[2374]*kernel[2]+tmp[2472]*kernel[3]+tmp[2473]*kernel[4]+tmp[2474]*kernel[5]+tmp[2572]*kernel[6]+tmp[2573]*kernel[7]+tmp[2574]*kernel[8];
				ans[2474]<=tmp[2373]*kernel[0]+tmp[2374]*kernel[1]+tmp[2375]*kernel[2]+tmp[2473]*kernel[3]+tmp[2474]*kernel[4]+tmp[2475]*kernel[5]+tmp[2573]*kernel[6]+tmp[2574]*kernel[7]+tmp[2575]*kernel[8];
				ans[2475]<=tmp[2374]*kernel[0]+tmp[2375]*kernel[1]+tmp[2376]*kernel[2]+tmp[2474]*kernel[3]+tmp[2475]*kernel[4]+tmp[2476]*kernel[5]+tmp[2574]*kernel[6]+tmp[2575]*kernel[7]+tmp[2576]*kernel[8];
				ans[2476]<=tmp[2375]*kernel[0]+tmp[2376]*kernel[1]+tmp[2377]*kernel[2]+tmp[2475]*kernel[3]+tmp[2476]*kernel[4]+tmp[2477]*kernel[5]+tmp[2575]*kernel[6]+tmp[2576]*kernel[7]+tmp[2577]*kernel[8];
				ans[2477]<=tmp[2376]*kernel[0]+tmp[2377]*kernel[1]+tmp[2378]*kernel[2]+tmp[2476]*kernel[3]+tmp[2477]*kernel[4]+tmp[2478]*kernel[5]+tmp[2576]*kernel[6]+tmp[2577]*kernel[7]+tmp[2578]*kernel[8];
				ans[2478]<=tmp[2377]*kernel[0]+tmp[2378]*kernel[1]+tmp[2379]*kernel[2]+tmp[2477]*kernel[3]+tmp[2478]*kernel[4]+tmp[2479]*kernel[5]+tmp[2577]*kernel[6]+tmp[2578]*kernel[7]+tmp[2579]*kernel[8];
				ans[2479]<=tmp[2378]*kernel[0]+tmp[2379]*kernel[1]+tmp[2380]*kernel[2]+tmp[2478]*kernel[3]+tmp[2479]*kernel[4]+tmp[2480]*kernel[5]+tmp[2578]*kernel[6]+tmp[2579]*kernel[7]+tmp[2580]*kernel[8];
				ans[2480]<=tmp[2379]*kernel[0]+tmp[2380]*kernel[1]+tmp[2381]*kernel[2]+tmp[2479]*kernel[3]+tmp[2480]*kernel[4]+tmp[2481]*kernel[5]+tmp[2579]*kernel[6]+tmp[2580]*kernel[7]+tmp[2581]*kernel[8];
				ans[2481]<=tmp[2380]*kernel[0]+tmp[2381]*kernel[1]+tmp[2382]*kernel[2]+tmp[2480]*kernel[3]+tmp[2481]*kernel[4]+tmp[2482]*kernel[5]+tmp[2580]*kernel[6]+tmp[2581]*kernel[7]+tmp[2582]*kernel[8];
				ans[2482]<=tmp[2381]*kernel[0]+tmp[2382]*kernel[1]+tmp[2383]*kernel[2]+tmp[2481]*kernel[3]+tmp[2482]*kernel[4]+tmp[2483]*kernel[5]+tmp[2581]*kernel[6]+tmp[2582]*kernel[7]+tmp[2583]*kernel[8];
				ans[2483]<=tmp[2382]*kernel[0]+tmp[2383]*kernel[1]+tmp[2384]*kernel[2]+tmp[2482]*kernel[3]+tmp[2483]*kernel[4]+tmp[2484]*kernel[5]+tmp[2582]*kernel[6]+tmp[2583]*kernel[7]+tmp[2584]*kernel[8];
				ans[2484]<=tmp[2383]*kernel[0]+tmp[2384]*kernel[1]+tmp[2385]*kernel[2]+tmp[2483]*kernel[3]+tmp[2484]*kernel[4]+tmp[2485]*kernel[5]+tmp[2583]*kernel[6]+tmp[2584]*kernel[7]+tmp[2585]*kernel[8];
				ans[2485]<=tmp[2384]*kernel[0]+tmp[2385]*kernel[1]+tmp[2386]*kernel[2]+tmp[2484]*kernel[3]+tmp[2485]*kernel[4]+tmp[2486]*kernel[5]+tmp[2584]*kernel[6]+tmp[2585]*kernel[7]+tmp[2586]*kernel[8];
				ans[2486]<=tmp[2385]*kernel[0]+tmp[2386]*kernel[1]+tmp[2387]*kernel[2]+tmp[2485]*kernel[3]+tmp[2486]*kernel[4]+tmp[2487]*kernel[5]+tmp[2585]*kernel[6]+tmp[2586]*kernel[7]+tmp[2587]*kernel[8];
				ans[2487]<=tmp[2386]*kernel[0]+tmp[2387]*kernel[1]+tmp[2388]*kernel[2]+tmp[2486]*kernel[3]+tmp[2487]*kernel[4]+tmp[2488]*kernel[5]+tmp[2586]*kernel[6]+tmp[2587]*kernel[7]+tmp[2588]*kernel[8];
				ans[2488]<=tmp[2387]*kernel[0]+tmp[2388]*kernel[1]+tmp[2389]*kernel[2]+tmp[2487]*kernel[3]+tmp[2488]*kernel[4]+tmp[2489]*kernel[5]+tmp[2587]*kernel[6]+tmp[2588]*kernel[7]+tmp[2589]*kernel[8];
				ans[2489]<=tmp[2388]*kernel[0]+tmp[2389]*kernel[1]+tmp[2390]*kernel[2]+tmp[2488]*kernel[3]+tmp[2489]*kernel[4]+tmp[2490]*kernel[5]+tmp[2588]*kernel[6]+tmp[2589]*kernel[7]+tmp[2590]*kernel[8];
				ans[2490]<=tmp[2389]*kernel[0]+tmp[2390]*kernel[1]+tmp[2391]*kernel[2]+tmp[2489]*kernel[3]+tmp[2490]*kernel[4]+tmp[2491]*kernel[5]+tmp[2589]*kernel[6]+tmp[2590]*kernel[7]+tmp[2591]*kernel[8];
				ans[2491]<=tmp[2390]*kernel[0]+tmp[2391]*kernel[1]+tmp[2392]*kernel[2]+tmp[2490]*kernel[3]+tmp[2491]*kernel[4]+tmp[2492]*kernel[5]+tmp[2590]*kernel[6]+tmp[2591]*kernel[7]+tmp[2592]*kernel[8];
				ans[2492]<=tmp[2391]*kernel[0]+tmp[2392]*kernel[1]+tmp[2393]*kernel[2]+tmp[2491]*kernel[3]+tmp[2492]*kernel[4]+tmp[2493]*kernel[5]+tmp[2591]*kernel[6]+tmp[2592]*kernel[7]+tmp[2593]*kernel[8];
				ans[2493]<=tmp[2392]*kernel[0]+tmp[2393]*kernel[1]+tmp[2394]*kernel[2]+tmp[2492]*kernel[3]+tmp[2493]*kernel[4]+tmp[2494]*kernel[5]+tmp[2592]*kernel[6]+tmp[2593]*kernel[7]+tmp[2594]*kernel[8];
				ans[2494]<=tmp[2393]*kernel[0]+tmp[2394]*kernel[1]+tmp[2395]*kernel[2]+tmp[2493]*kernel[3]+tmp[2494]*kernel[4]+tmp[2495]*kernel[5]+tmp[2593]*kernel[6]+tmp[2594]*kernel[7]+tmp[2595]*kernel[8];
				ans[2495]<=tmp[2394]*kernel[0]+tmp[2395]*kernel[1]+tmp[2396]*kernel[2]+tmp[2494]*kernel[3]+tmp[2495]*kernel[4]+tmp[2496]*kernel[5]+tmp[2594]*kernel[6]+tmp[2595]*kernel[7]+tmp[2596]*kernel[8];
				ans[2496]<=tmp[2395]*kernel[0]+tmp[2396]*kernel[1]+tmp[2397]*kernel[2]+tmp[2495]*kernel[3]+tmp[2496]*kernel[4]+tmp[2497]*kernel[5]+tmp[2595]*kernel[6]+tmp[2596]*kernel[7]+tmp[2597]*kernel[8];
				ans[2497]<=tmp[2396]*kernel[0]+tmp[2397]*kernel[1]+tmp[2398]*kernel[2]+tmp[2496]*kernel[3]+tmp[2497]*kernel[4]+tmp[2498]*kernel[5]+tmp[2596]*kernel[6]+tmp[2597]*kernel[7]+tmp[2598]*kernel[8];
				ans[2498]<=tmp[2397]*kernel[0]+tmp[2398]*kernel[1]+tmp[2399]*kernel[2]+tmp[2497]*kernel[3]+tmp[2498]*kernel[4]+tmp[2499]*kernel[5]+tmp[2597]*kernel[6]+tmp[2598]*kernel[7]+tmp[2599]*kernel[8];
				ans[2499]<=tmp[2398]*kernel[0]+tmp[2399]*kernel[1]+tmp[2498]*kernel[3]+tmp[2499]*kernel[4]+tmp[2598]*kernel[6]+tmp[2599]*kernel[7];
				ans[2500]<=tmp[2400]*kernel[1]+tmp[2401]*kernel[2]+tmp[2500]*kernel[4]+tmp[2501]*kernel[5]+tmp[2600]*kernel[7]+tmp[2601]*kernel[8];
				ans[2501]<=tmp[2400]*kernel[0]+tmp[2401]*kernel[1]+tmp[2402]*kernel[2]+tmp[2500]*kernel[3]+tmp[2501]*kernel[4]+tmp[2502]*kernel[5]+tmp[2600]*kernel[6]+tmp[2601]*kernel[7]+tmp[2602]*kernel[8];
				ans[2502]<=tmp[2401]*kernel[0]+tmp[2402]*kernel[1]+tmp[2403]*kernel[2]+tmp[2501]*kernel[3]+tmp[2502]*kernel[4]+tmp[2503]*kernel[5]+tmp[2601]*kernel[6]+tmp[2602]*kernel[7]+tmp[2603]*kernel[8];
				ans[2503]<=tmp[2402]*kernel[0]+tmp[2403]*kernel[1]+tmp[2404]*kernel[2]+tmp[2502]*kernel[3]+tmp[2503]*kernel[4]+tmp[2504]*kernel[5]+tmp[2602]*kernel[6]+tmp[2603]*kernel[7]+tmp[2604]*kernel[8];
				ans[2504]<=tmp[2403]*kernel[0]+tmp[2404]*kernel[1]+tmp[2405]*kernel[2]+tmp[2503]*kernel[3]+tmp[2504]*kernel[4]+tmp[2505]*kernel[5]+tmp[2603]*kernel[6]+tmp[2604]*kernel[7]+tmp[2605]*kernel[8];
				ans[2505]<=tmp[2404]*kernel[0]+tmp[2405]*kernel[1]+tmp[2406]*kernel[2]+tmp[2504]*kernel[3]+tmp[2505]*kernel[4]+tmp[2506]*kernel[5]+tmp[2604]*kernel[6]+tmp[2605]*kernel[7]+tmp[2606]*kernel[8];
				ans[2506]<=tmp[2405]*kernel[0]+tmp[2406]*kernel[1]+tmp[2407]*kernel[2]+tmp[2505]*kernel[3]+tmp[2506]*kernel[4]+tmp[2507]*kernel[5]+tmp[2605]*kernel[6]+tmp[2606]*kernel[7]+tmp[2607]*kernel[8];
				ans[2507]<=tmp[2406]*kernel[0]+tmp[2407]*kernel[1]+tmp[2408]*kernel[2]+tmp[2506]*kernel[3]+tmp[2507]*kernel[4]+tmp[2508]*kernel[5]+tmp[2606]*kernel[6]+tmp[2607]*kernel[7]+tmp[2608]*kernel[8];
				ans[2508]<=tmp[2407]*kernel[0]+tmp[2408]*kernel[1]+tmp[2409]*kernel[2]+tmp[2507]*kernel[3]+tmp[2508]*kernel[4]+tmp[2509]*kernel[5]+tmp[2607]*kernel[6]+tmp[2608]*kernel[7]+tmp[2609]*kernel[8];
				ans[2509]<=tmp[2408]*kernel[0]+tmp[2409]*kernel[1]+tmp[2410]*kernel[2]+tmp[2508]*kernel[3]+tmp[2509]*kernel[4]+tmp[2510]*kernel[5]+tmp[2608]*kernel[6]+tmp[2609]*kernel[7]+tmp[2610]*kernel[8];
				ans[2510]<=tmp[2409]*kernel[0]+tmp[2410]*kernel[1]+tmp[2411]*kernel[2]+tmp[2509]*kernel[3]+tmp[2510]*kernel[4]+tmp[2511]*kernel[5]+tmp[2609]*kernel[6]+tmp[2610]*kernel[7]+tmp[2611]*kernel[8];
				ans[2511]<=tmp[2410]*kernel[0]+tmp[2411]*kernel[1]+tmp[2412]*kernel[2]+tmp[2510]*kernel[3]+tmp[2511]*kernel[4]+tmp[2512]*kernel[5]+tmp[2610]*kernel[6]+tmp[2611]*kernel[7]+tmp[2612]*kernel[8];
				ans[2512]<=tmp[2411]*kernel[0]+tmp[2412]*kernel[1]+tmp[2413]*kernel[2]+tmp[2511]*kernel[3]+tmp[2512]*kernel[4]+tmp[2513]*kernel[5]+tmp[2611]*kernel[6]+tmp[2612]*kernel[7]+tmp[2613]*kernel[8];
				ans[2513]<=tmp[2412]*kernel[0]+tmp[2413]*kernel[1]+tmp[2414]*kernel[2]+tmp[2512]*kernel[3]+tmp[2513]*kernel[4]+tmp[2514]*kernel[5]+tmp[2612]*kernel[6]+tmp[2613]*kernel[7]+tmp[2614]*kernel[8];
				ans[2514]<=tmp[2413]*kernel[0]+tmp[2414]*kernel[1]+tmp[2415]*kernel[2]+tmp[2513]*kernel[3]+tmp[2514]*kernel[4]+tmp[2515]*kernel[5]+tmp[2613]*kernel[6]+tmp[2614]*kernel[7]+tmp[2615]*kernel[8];
				ans[2515]<=tmp[2414]*kernel[0]+tmp[2415]*kernel[1]+tmp[2416]*kernel[2]+tmp[2514]*kernel[3]+tmp[2515]*kernel[4]+tmp[2516]*kernel[5]+tmp[2614]*kernel[6]+tmp[2615]*kernel[7]+tmp[2616]*kernel[8];
				ans[2516]<=tmp[2415]*kernel[0]+tmp[2416]*kernel[1]+tmp[2417]*kernel[2]+tmp[2515]*kernel[3]+tmp[2516]*kernel[4]+tmp[2517]*kernel[5]+tmp[2615]*kernel[6]+tmp[2616]*kernel[7]+tmp[2617]*kernel[8];
				ans[2517]<=tmp[2416]*kernel[0]+tmp[2417]*kernel[1]+tmp[2418]*kernel[2]+tmp[2516]*kernel[3]+tmp[2517]*kernel[4]+tmp[2518]*kernel[5]+tmp[2616]*kernel[6]+tmp[2617]*kernel[7]+tmp[2618]*kernel[8];
				ans[2518]<=tmp[2417]*kernel[0]+tmp[2418]*kernel[1]+tmp[2419]*kernel[2]+tmp[2517]*kernel[3]+tmp[2518]*kernel[4]+tmp[2519]*kernel[5]+tmp[2617]*kernel[6]+tmp[2618]*kernel[7]+tmp[2619]*kernel[8];
				ans[2519]<=tmp[2418]*kernel[0]+tmp[2419]*kernel[1]+tmp[2420]*kernel[2]+tmp[2518]*kernel[3]+tmp[2519]*kernel[4]+tmp[2520]*kernel[5]+tmp[2618]*kernel[6]+tmp[2619]*kernel[7]+tmp[2620]*kernel[8];
				ans[2520]<=tmp[2419]*kernel[0]+tmp[2420]*kernel[1]+tmp[2421]*kernel[2]+tmp[2519]*kernel[3]+tmp[2520]*kernel[4]+tmp[2521]*kernel[5]+tmp[2619]*kernel[6]+tmp[2620]*kernel[7]+tmp[2621]*kernel[8];
				ans[2521]<=tmp[2420]*kernel[0]+tmp[2421]*kernel[1]+tmp[2422]*kernel[2]+tmp[2520]*kernel[3]+tmp[2521]*kernel[4]+tmp[2522]*kernel[5]+tmp[2620]*kernel[6]+tmp[2621]*kernel[7]+tmp[2622]*kernel[8];
				ans[2522]<=tmp[2421]*kernel[0]+tmp[2422]*kernel[1]+tmp[2423]*kernel[2]+tmp[2521]*kernel[3]+tmp[2522]*kernel[4]+tmp[2523]*kernel[5]+tmp[2621]*kernel[6]+tmp[2622]*kernel[7]+tmp[2623]*kernel[8];
				ans[2523]<=tmp[2422]*kernel[0]+tmp[2423]*kernel[1]+tmp[2424]*kernel[2]+tmp[2522]*kernel[3]+tmp[2523]*kernel[4]+tmp[2524]*kernel[5]+tmp[2622]*kernel[6]+tmp[2623]*kernel[7]+tmp[2624]*kernel[8];
				ans[2524]<=tmp[2423]*kernel[0]+tmp[2424]*kernel[1]+tmp[2425]*kernel[2]+tmp[2523]*kernel[3]+tmp[2524]*kernel[4]+tmp[2525]*kernel[5]+tmp[2623]*kernel[6]+tmp[2624]*kernel[7]+tmp[2625]*kernel[8];
				ans[2525]<=tmp[2424]*kernel[0]+tmp[2425]*kernel[1]+tmp[2426]*kernel[2]+tmp[2524]*kernel[3]+tmp[2525]*kernel[4]+tmp[2526]*kernel[5]+tmp[2624]*kernel[6]+tmp[2625]*kernel[7]+tmp[2626]*kernel[8];
				ans[2526]<=tmp[2425]*kernel[0]+tmp[2426]*kernel[1]+tmp[2427]*kernel[2]+tmp[2525]*kernel[3]+tmp[2526]*kernel[4]+tmp[2527]*kernel[5]+tmp[2625]*kernel[6]+tmp[2626]*kernel[7]+tmp[2627]*kernel[8];
				ans[2527]<=tmp[2426]*kernel[0]+tmp[2427]*kernel[1]+tmp[2428]*kernel[2]+tmp[2526]*kernel[3]+tmp[2527]*kernel[4]+tmp[2528]*kernel[5]+tmp[2626]*kernel[6]+tmp[2627]*kernel[7]+tmp[2628]*kernel[8];
				ans[2528]<=tmp[2427]*kernel[0]+tmp[2428]*kernel[1]+tmp[2429]*kernel[2]+tmp[2527]*kernel[3]+tmp[2528]*kernel[4]+tmp[2529]*kernel[5]+tmp[2627]*kernel[6]+tmp[2628]*kernel[7]+tmp[2629]*kernel[8];
				ans[2529]<=tmp[2428]*kernel[0]+tmp[2429]*kernel[1]+tmp[2430]*kernel[2]+tmp[2528]*kernel[3]+tmp[2529]*kernel[4]+tmp[2530]*kernel[5]+tmp[2628]*kernel[6]+tmp[2629]*kernel[7]+tmp[2630]*kernel[8];
				ans[2530]<=tmp[2429]*kernel[0]+tmp[2430]*kernel[1]+tmp[2431]*kernel[2]+tmp[2529]*kernel[3]+tmp[2530]*kernel[4]+tmp[2531]*kernel[5]+tmp[2629]*kernel[6]+tmp[2630]*kernel[7]+tmp[2631]*kernel[8];
				ans[2531]<=tmp[2430]*kernel[0]+tmp[2431]*kernel[1]+tmp[2432]*kernel[2]+tmp[2530]*kernel[3]+tmp[2531]*kernel[4]+tmp[2532]*kernel[5]+tmp[2630]*kernel[6]+tmp[2631]*kernel[7]+tmp[2632]*kernel[8];
				ans[2532]<=tmp[2431]*kernel[0]+tmp[2432]*kernel[1]+tmp[2433]*kernel[2]+tmp[2531]*kernel[3]+tmp[2532]*kernel[4]+tmp[2533]*kernel[5]+tmp[2631]*kernel[6]+tmp[2632]*kernel[7]+tmp[2633]*kernel[8];
				ans[2533]<=tmp[2432]*kernel[0]+tmp[2433]*kernel[1]+tmp[2434]*kernel[2]+tmp[2532]*kernel[3]+tmp[2533]*kernel[4]+tmp[2534]*kernel[5]+tmp[2632]*kernel[6]+tmp[2633]*kernel[7]+tmp[2634]*kernel[8];
				ans[2534]<=tmp[2433]*kernel[0]+tmp[2434]*kernel[1]+tmp[2435]*kernel[2]+tmp[2533]*kernel[3]+tmp[2534]*kernel[4]+tmp[2535]*kernel[5]+tmp[2633]*kernel[6]+tmp[2634]*kernel[7]+tmp[2635]*kernel[8];
				ans[2535]<=tmp[2434]*kernel[0]+tmp[2435]*kernel[1]+tmp[2436]*kernel[2]+tmp[2534]*kernel[3]+tmp[2535]*kernel[4]+tmp[2536]*kernel[5]+tmp[2634]*kernel[6]+tmp[2635]*kernel[7]+tmp[2636]*kernel[8];
				ans[2536]<=tmp[2435]*kernel[0]+tmp[2436]*kernel[1]+tmp[2437]*kernel[2]+tmp[2535]*kernel[3]+tmp[2536]*kernel[4]+tmp[2537]*kernel[5]+tmp[2635]*kernel[6]+tmp[2636]*kernel[7]+tmp[2637]*kernel[8];
				ans[2537]<=tmp[2436]*kernel[0]+tmp[2437]*kernel[1]+tmp[2438]*kernel[2]+tmp[2536]*kernel[3]+tmp[2537]*kernel[4]+tmp[2538]*kernel[5]+tmp[2636]*kernel[6]+tmp[2637]*kernel[7]+tmp[2638]*kernel[8];
				ans[2538]<=tmp[2437]*kernel[0]+tmp[2438]*kernel[1]+tmp[2439]*kernel[2]+tmp[2537]*kernel[3]+tmp[2538]*kernel[4]+tmp[2539]*kernel[5]+tmp[2637]*kernel[6]+tmp[2638]*kernel[7]+tmp[2639]*kernel[8];
				ans[2539]<=tmp[2438]*kernel[0]+tmp[2439]*kernel[1]+tmp[2440]*kernel[2]+tmp[2538]*kernel[3]+tmp[2539]*kernel[4]+tmp[2540]*kernel[5]+tmp[2638]*kernel[6]+tmp[2639]*kernel[7]+tmp[2640]*kernel[8];
				ans[2540]<=tmp[2439]*kernel[0]+tmp[2440]*kernel[1]+tmp[2441]*kernel[2]+tmp[2539]*kernel[3]+tmp[2540]*kernel[4]+tmp[2541]*kernel[5]+tmp[2639]*kernel[6]+tmp[2640]*kernel[7]+tmp[2641]*kernel[8];
				ans[2541]<=tmp[2440]*kernel[0]+tmp[2441]*kernel[1]+tmp[2442]*kernel[2]+tmp[2540]*kernel[3]+tmp[2541]*kernel[4]+tmp[2542]*kernel[5]+tmp[2640]*kernel[6]+tmp[2641]*kernel[7]+tmp[2642]*kernel[8];
				ans[2542]<=tmp[2441]*kernel[0]+tmp[2442]*kernel[1]+tmp[2443]*kernel[2]+tmp[2541]*kernel[3]+tmp[2542]*kernel[4]+tmp[2543]*kernel[5]+tmp[2641]*kernel[6]+tmp[2642]*kernel[7]+tmp[2643]*kernel[8];
				ans[2543]<=tmp[2442]*kernel[0]+tmp[2443]*kernel[1]+tmp[2444]*kernel[2]+tmp[2542]*kernel[3]+tmp[2543]*kernel[4]+tmp[2544]*kernel[5]+tmp[2642]*kernel[6]+tmp[2643]*kernel[7]+tmp[2644]*kernel[8];
				ans[2544]<=tmp[2443]*kernel[0]+tmp[2444]*kernel[1]+tmp[2445]*kernel[2]+tmp[2543]*kernel[3]+tmp[2544]*kernel[4]+tmp[2545]*kernel[5]+tmp[2643]*kernel[6]+tmp[2644]*kernel[7]+tmp[2645]*kernel[8];
				ans[2545]<=tmp[2444]*kernel[0]+tmp[2445]*kernel[1]+tmp[2446]*kernel[2]+tmp[2544]*kernel[3]+tmp[2545]*kernel[4]+tmp[2546]*kernel[5]+tmp[2644]*kernel[6]+tmp[2645]*kernel[7]+tmp[2646]*kernel[8];
				ans[2546]<=tmp[2445]*kernel[0]+tmp[2446]*kernel[1]+tmp[2447]*kernel[2]+tmp[2545]*kernel[3]+tmp[2546]*kernel[4]+tmp[2547]*kernel[5]+tmp[2645]*kernel[6]+tmp[2646]*kernel[7]+tmp[2647]*kernel[8];
				ans[2547]<=tmp[2446]*kernel[0]+tmp[2447]*kernel[1]+tmp[2448]*kernel[2]+tmp[2546]*kernel[3]+tmp[2547]*kernel[4]+tmp[2548]*kernel[5]+tmp[2646]*kernel[6]+tmp[2647]*kernel[7]+tmp[2648]*kernel[8];
				ans[2548]<=tmp[2447]*kernel[0]+tmp[2448]*kernel[1]+tmp[2449]*kernel[2]+tmp[2547]*kernel[3]+tmp[2548]*kernel[4]+tmp[2549]*kernel[5]+tmp[2647]*kernel[6]+tmp[2648]*kernel[7]+tmp[2649]*kernel[8];
				ans[2549]<=tmp[2448]*kernel[0]+tmp[2449]*kernel[1]+tmp[2450]*kernel[2]+tmp[2548]*kernel[3]+tmp[2549]*kernel[4]+tmp[2550]*kernel[5]+tmp[2648]*kernel[6]+tmp[2649]*kernel[7]+tmp[2650]*kernel[8];
				ans[2550]<=tmp[2449]*kernel[0]+tmp[2450]*kernel[1]+tmp[2451]*kernel[2]+tmp[2549]*kernel[3]+tmp[2550]*kernel[4]+tmp[2551]*kernel[5]+tmp[2649]*kernel[6]+tmp[2650]*kernel[7]+tmp[2651]*kernel[8];
				ans[2551]<=tmp[2450]*kernel[0]+tmp[2451]*kernel[1]+tmp[2452]*kernel[2]+tmp[2550]*kernel[3]+tmp[2551]*kernel[4]+tmp[2552]*kernel[5]+tmp[2650]*kernel[6]+tmp[2651]*kernel[7]+tmp[2652]*kernel[8];
				ans[2552]<=tmp[2451]*kernel[0]+tmp[2452]*kernel[1]+tmp[2453]*kernel[2]+tmp[2551]*kernel[3]+tmp[2552]*kernel[4]+tmp[2553]*kernel[5]+tmp[2651]*kernel[6]+tmp[2652]*kernel[7]+tmp[2653]*kernel[8];
				ans[2553]<=tmp[2452]*kernel[0]+tmp[2453]*kernel[1]+tmp[2454]*kernel[2]+tmp[2552]*kernel[3]+tmp[2553]*kernel[4]+tmp[2554]*kernel[5]+tmp[2652]*kernel[6]+tmp[2653]*kernel[7]+tmp[2654]*kernel[8];
				ans[2554]<=tmp[2453]*kernel[0]+tmp[2454]*kernel[1]+tmp[2455]*kernel[2]+tmp[2553]*kernel[3]+tmp[2554]*kernel[4]+tmp[2555]*kernel[5]+tmp[2653]*kernel[6]+tmp[2654]*kernel[7]+tmp[2655]*kernel[8];
				ans[2555]<=tmp[2454]*kernel[0]+tmp[2455]*kernel[1]+tmp[2456]*kernel[2]+tmp[2554]*kernel[3]+tmp[2555]*kernel[4]+tmp[2556]*kernel[5]+tmp[2654]*kernel[6]+tmp[2655]*kernel[7]+tmp[2656]*kernel[8];
				ans[2556]<=tmp[2455]*kernel[0]+tmp[2456]*kernel[1]+tmp[2457]*kernel[2]+tmp[2555]*kernel[3]+tmp[2556]*kernel[4]+tmp[2557]*kernel[5]+tmp[2655]*kernel[6]+tmp[2656]*kernel[7]+tmp[2657]*kernel[8];
				ans[2557]<=tmp[2456]*kernel[0]+tmp[2457]*kernel[1]+tmp[2458]*kernel[2]+tmp[2556]*kernel[3]+tmp[2557]*kernel[4]+tmp[2558]*kernel[5]+tmp[2656]*kernel[6]+tmp[2657]*kernel[7]+tmp[2658]*kernel[8];
				ans[2558]<=tmp[2457]*kernel[0]+tmp[2458]*kernel[1]+tmp[2459]*kernel[2]+tmp[2557]*kernel[3]+tmp[2558]*kernel[4]+tmp[2559]*kernel[5]+tmp[2657]*kernel[6]+tmp[2658]*kernel[7]+tmp[2659]*kernel[8];
				ans[2559]<=tmp[2458]*kernel[0]+tmp[2459]*kernel[1]+tmp[2460]*kernel[2]+tmp[2558]*kernel[3]+tmp[2559]*kernel[4]+tmp[2560]*kernel[5]+tmp[2658]*kernel[6]+tmp[2659]*kernel[7]+tmp[2660]*kernel[8];
				ans[2560]<=tmp[2459]*kernel[0]+tmp[2460]*kernel[1]+tmp[2461]*kernel[2]+tmp[2559]*kernel[3]+tmp[2560]*kernel[4]+tmp[2561]*kernel[5]+tmp[2659]*kernel[6]+tmp[2660]*kernel[7]+tmp[2661]*kernel[8];
				ans[2561]<=tmp[2460]*kernel[0]+tmp[2461]*kernel[1]+tmp[2462]*kernel[2]+tmp[2560]*kernel[3]+tmp[2561]*kernel[4]+tmp[2562]*kernel[5]+tmp[2660]*kernel[6]+tmp[2661]*kernel[7]+tmp[2662]*kernel[8];
				ans[2562]<=tmp[2461]*kernel[0]+tmp[2462]*kernel[1]+tmp[2463]*kernel[2]+tmp[2561]*kernel[3]+tmp[2562]*kernel[4]+tmp[2563]*kernel[5]+tmp[2661]*kernel[6]+tmp[2662]*kernel[7]+tmp[2663]*kernel[8];
				ans[2563]<=tmp[2462]*kernel[0]+tmp[2463]*kernel[1]+tmp[2464]*kernel[2]+tmp[2562]*kernel[3]+tmp[2563]*kernel[4]+tmp[2564]*kernel[5]+tmp[2662]*kernel[6]+tmp[2663]*kernel[7]+tmp[2664]*kernel[8];
				ans[2564]<=tmp[2463]*kernel[0]+tmp[2464]*kernel[1]+tmp[2465]*kernel[2]+tmp[2563]*kernel[3]+tmp[2564]*kernel[4]+tmp[2565]*kernel[5]+tmp[2663]*kernel[6]+tmp[2664]*kernel[7]+tmp[2665]*kernel[8];
				ans[2565]<=tmp[2464]*kernel[0]+tmp[2465]*kernel[1]+tmp[2466]*kernel[2]+tmp[2564]*kernel[3]+tmp[2565]*kernel[4]+tmp[2566]*kernel[5]+tmp[2664]*kernel[6]+tmp[2665]*kernel[7]+tmp[2666]*kernel[8];
				ans[2566]<=tmp[2465]*kernel[0]+tmp[2466]*kernel[1]+tmp[2467]*kernel[2]+tmp[2565]*kernel[3]+tmp[2566]*kernel[4]+tmp[2567]*kernel[5]+tmp[2665]*kernel[6]+tmp[2666]*kernel[7]+tmp[2667]*kernel[8];
				ans[2567]<=tmp[2466]*kernel[0]+tmp[2467]*kernel[1]+tmp[2468]*kernel[2]+tmp[2566]*kernel[3]+tmp[2567]*kernel[4]+tmp[2568]*kernel[5]+tmp[2666]*kernel[6]+tmp[2667]*kernel[7]+tmp[2668]*kernel[8];
				ans[2568]<=tmp[2467]*kernel[0]+tmp[2468]*kernel[1]+tmp[2469]*kernel[2]+tmp[2567]*kernel[3]+tmp[2568]*kernel[4]+tmp[2569]*kernel[5]+tmp[2667]*kernel[6]+tmp[2668]*kernel[7]+tmp[2669]*kernel[8];
				ans[2569]<=tmp[2468]*kernel[0]+tmp[2469]*kernel[1]+tmp[2470]*kernel[2]+tmp[2568]*kernel[3]+tmp[2569]*kernel[4]+tmp[2570]*kernel[5]+tmp[2668]*kernel[6]+tmp[2669]*kernel[7]+tmp[2670]*kernel[8];
				ans[2570]<=tmp[2469]*kernel[0]+tmp[2470]*kernel[1]+tmp[2471]*kernel[2]+tmp[2569]*kernel[3]+tmp[2570]*kernel[4]+tmp[2571]*kernel[5]+tmp[2669]*kernel[6]+tmp[2670]*kernel[7]+tmp[2671]*kernel[8];
				ans[2571]<=tmp[2470]*kernel[0]+tmp[2471]*kernel[1]+tmp[2472]*kernel[2]+tmp[2570]*kernel[3]+tmp[2571]*kernel[4]+tmp[2572]*kernel[5]+tmp[2670]*kernel[6]+tmp[2671]*kernel[7]+tmp[2672]*kernel[8];
				ans[2572]<=tmp[2471]*kernel[0]+tmp[2472]*kernel[1]+tmp[2473]*kernel[2]+tmp[2571]*kernel[3]+tmp[2572]*kernel[4]+tmp[2573]*kernel[5]+tmp[2671]*kernel[6]+tmp[2672]*kernel[7]+tmp[2673]*kernel[8];
				ans[2573]<=tmp[2472]*kernel[0]+tmp[2473]*kernel[1]+tmp[2474]*kernel[2]+tmp[2572]*kernel[3]+tmp[2573]*kernel[4]+tmp[2574]*kernel[5]+tmp[2672]*kernel[6]+tmp[2673]*kernel[7]+tmp[2674]*kernel[8];
				ans[2574]<=tmp[2473]*kernel[0]+tmp[2474]*kernel[1]+tmp[2475]*kernel[2]+tmp[2573]*kernel[3]+tmp[2574]*kernel[4]+tmp[2575]*kernel[5]+tmp[2673]*kernel[6]+tmp[2674]*kernel[7]+tmp[2675]*kernel[8];
				ans[2575]<=tmp[2474]*kernel[0]+tmp[2475]*kernel[1]+tmp[2476]*kernel[2]+tmp[2574]*kernel[3]+tmp[2575]*kernel[4]+tmp[2576]*kernel[5]+tmp[2674]*kernel[6]+tmp[2675]*kernel[7]+tmp[2676]*kernel[8];
				ans[2576]<=tmp[2475]*kernel[0]+tmp[2476]*kernel[1]+tmp[2477]*kernel[2]+tmp[2575]*kernel[3]+tmp[2576]*kernel[4]+tmp[2577]*kernel[5]+tmp[2675]*kernel[6]+tmp[2676]*kernel[7]+tmp[2677]*kernel[8];
				ans[2577]<=tmp[2476]*kernel[0]+tmp[2477]*kernel[1]+tmp[2478]*kernel[2]+tmp[2576]*kernel[3]+tmp[2577]*kernel[4]+tmp[2578]*kernel[5]+tmp[2676]*kernel[6]+tmp[2677]*kernel[7]+tmp[2678]*kernel[8];
				ans[2578]<=tmp[2477]*kernel[0]+tmp[2478]*kernel[1]+tmp[2479]*kernel[2]+tmp[2577]*kernel[3]+tmp[2578]*kernel[4]+tmp[2579]*kernel[5]+tmp[2677]*kernel[6]+tmp[2678]*kernel[7]+tmp[2679]*kernel[8];
				ans[2579]<=tmp[2478]*kernel[0]+tmp[2479]*kernel[1]+tmp[2480]*kernel[2]+tmp[2578]*kernel[3]+tmp[2579]*kernel[4]+tmp[2580]*kernel[5]+tmp[2678]*kernel[6]+tmp[2679]*kernel[7]+tmp[2680]*kernel[8];
				ans[2580]<=tmp[2479]*kernel[0]+tmp[2480]*kernel[1]+tmp[2481]*kernel[2]+tmp[2579]*kernel[3]+tmp[2580]*kernel[4]+tmp[2581]*kernel[5]+tmp[2679]*kernel[6]+tmp[2680]*kernel[7]+tmp[2681]*kernel[8];
				ans[2581]<=tmp[2480]*kernel[0]+tmp[2481]*kernel[1]+tmp[2482]*kernel[2]+tmp[2580]*kernel[3]+tmp[2581]*kernel[4]+tmp[2582]*kernel[5]+tmp[2680]*kernel[6]+tmp[2681]*kernel[7]+tmp[2682]*kernel[8];
				ans[2582]<=tmp[2481]*kernel[0]+tmp[2482]*kernel[1]+tmp[2483]*kernel[2]+tmp[2581]*kernel[3]+tmp[2582]*kernel[4]+tmp[2583]*kernel[5]+tmp[2681]*kernel[6]+tmp[2682]*kernel[7]+tmp[2683]*kernel[8];
				ans[2583]<=tmp[2482]*kernel[0]+tmp[2483]*kernel[1]+tmp[2484]*kernel[2]+tmp[2582]*kernel[3]+tmp[2583]*kernel[4]+tmp[2584]*kernel[5]+tmp[2682]*kernel[6]+tmp[2683]*kernel[7]+tmp[2684]*kernel[8];
				ans[2584]<=tmp[2483]*kernel[0]+tmp[2484]*kernel[1]+tmp[2485]*kernel[2]+tmp[2583]*kernel[3]+tmp[2584]*kernel[4]+tmp[2585]*kernel[5]+tmp[2683]*kernel[6]+tmp[2684]*kernel[7]+tmp[2685]*kernel[8];
				ans[2585]<=tmp[2484]*kernel[0]+tmp[2485]*kernel[1]+tmp[2486]*kernel[2]+tmp[2584]*kernel[3]+tmp[2585]*kernel[4]+tmp[2586]*kernel[5]+tmp[2684]*kernel[6]+tmp[2685]*kernel[7]+tmp[2686]*kernel[8];
				ans[2586]<=tmp[2485]*kernel[0]+tmp[2486]*kernel[1]+tmp[2487]*kernel[2]+tmp[2585]*kernel[3]+tmp[2586]*kernel[4]+tmp[2587]*kernel[5]+tmp[2685]*kernel[6]+tmp[2686]*kernel[7]+tmp[2687]*kernel[8];
				ans[2587]<=tmp[2486]*kernel[0]+tmp[2487]*kernel[1]+tmp[2488]*kernel[2]+tmp[2586]*kernel[3]+tmp[2587]*kernel[4]+tmp[2588]*kernel[5]+tmp[2686]*kernel[6]+tmp[2687]*kernel[7]+tmp[2688]*kernel[8];
				ans[2588]<=tmp[2487]*kernel[0]+tmp[2488]*kernel[1]+tmp[2489]*kernel[2]+tmp[2587]*kernel[3]+tmp[2588]*kernel[4]+tmp[2589]*kernel[5]+tmp[2687]*kernel[6]+tmp[2688]*kernel[7]+tmp[2689]*kernel[8];
				ans[2589]<=tmp[2488]*kernel[0]+tmp[2489]*kernel[1]+tmp[2490]*kernel[2]+tmp[2588]*kernel[3]+tmp[2589]*kernel[4]+tmp[2590]*kernel[5]+tmp[2688]*kernel[6]+tmp[2689]*kernel[7]+tmp[2690]*kernel[8];
				ans[2590]<=tmp[2489]*kernel[0]+tmp[2490]*kernel[1]+tmp[2491]*kernel[2]+tmp[2589]*kernel[3]+tmp[2590]*kernel[4]+tmp[2591]*kernel[5]+tmp[2689]*kernel[6]+tmp[2690]*kernel[7]+tmp[2691]*kernel[8];
				ans[2591]<=tmp[2490]*kernel[0]+tmp[2491]*kernel[1]+tmp[2492]*kernel[2]+tmp[2590]*kernel[3]+tmp[2591]*kernel[4]+tmp[2592]*kernel[5]+tmp[2690]*kernel[6]+tmp[2691]*kernel[7]+tmp[2692]*kernel[8];
				ans[2592]<=tmp[2491]*kernel[0]+tmp[2492]*kernel[1]+tmp[2493]*kernel[2]+tmp[2591]*kernel[3]+tmp[2592]*kernel[4]+tmp[2593]*kernel[5]+tmp[2691]*kernel[6]+tmp[2692]*kernel[7]+tmp[2693]*kernel[8];
				ans[2593]<=tmp[2492]*kernel[0]+tmp[2493]*kernel[1]+tmp[2494]*kernel[2]+tmp[2592]*kernel[3]+tmp[2593]*kernel[4]+tmp[2594]*kernel[5]+tmp[2692]*kernel[6]+tmp[2693]*kernel[7]+tmp[2694]*kernel[8];
				ans[2594]<=tmp[2493]*kernel[0]+tmp[2494]*kernel[1]+tmp[2495]*kernel[2]+tmp[2593]*kernel[3]+tmp[2594]*kernel[4]+tmp[2595]*kernel[5]+tmp[2693]*kernel[6]+tmp[2694]*kernel[7]+tmp[2695]*kernel[8];
				ans[2595]<=tmp[2494]*kernel[0]+tmp[2495]*kernel[1]+tmp[2496]*kernel[2]+tmp[2594]*kernel[3]+tmp[2595]*kernel[4]+tmp[2596]*kernel[5]+tmp[2694]*kernel[6]+tmp[2695]*kernel[7]+tmp[2696]*kernel[8];
				ans[2596]<=tmp[2495]*kernel[0]+tmp[2496]*kernel[1]+tmp[2497]*kernel[2]+tmp[2595]*kernel[3]+tmp[2596]*kernel[4]+tmp[2597]*kernel[5]+tmp[2695]*kernel[6]+tmp[2696]*kernel[7]+tmp[2697]*kernel[8];
				ans[2597]<=tmp[2496]*kernel[0]+tmp[2497]*kernel[1]+tmp[2498]*kernel[2]+tmp[2596]*kernel[3]+tmp[2597]*kernel[4]+tmp[2598]*kernel[5]+tmp[2696]*kernel[6]+tmp[2697]*kernel[7]+tmp[2698]*kernel[8];
				ans[2598]<=tmp[2497]*kernel[0]+tmp[2498]*kernel[1]+tmp[2499]*kernel[2]+tmp[2597]*kernel[3]+tmp[2598]*kernel[4]+tmp[2599]*kernel[5]+tmp[2697]*kernel[6]+tmp[2698]*kernel[7]+tmp[2699]*kernel[8];
				ans[2599]<=tmp[2498]*kernel[0]+tmp[2499]*kernel[1]+tmp[2598]*kernel[3]+tmp[2599]*kernel[4]+tmp[2698]*kernel[6]+tmp[2699]*kernel[7];
				ans[2600]<=tmp[2500]*kernel[1]+tmp[2501]*kernel[2]+tmp[2600]*kernel[4]+tmp[2601]*kernel[5]+tmp[2700]*kernel[7]+tmp[2701]*kernel[8];
				ans[2601]<=tmp[2500]*kernel[0]+tmp[2501]*kernel[1]+tmp[2502]*kernel[2]+tmp[2600]*kernel[3]+tmp[2601]*kernel[4]+tmp[2602]*kernel[5]+tmp[2700]*kernel[6]+tmp[2701]*kernel[7]+tmp[2702]*kernel[8];
				ans[2602]<=tmp[2501]*kernel[0]+tmp[2502]*kernel[1]+tmp[2503]*kernel[2]+tmp[2601]*kernel[3]+tmp[2602]*kernel[4]+tmp[2603]*kernel[5]+tmp[2701]*kernel[6]+tmp[2702]*kernel[7]+tmp[2703]*kernel[8];
				ans[2603]<=tmp[2502]*kernel[0]+tmp[2503]*kernel[1]+tmp[2504]*kernel[2]+tmp[2602]*kernel[3]+tmp[2603]*kernel[4]+tmp[2604]*kernel[5]+tmp[2702]*kernel[6]+tmp[2703]*kernel[7]+tmp[2704]*kernel[8];
				ans[2604]<=tmp[2503]*kernel[0]+tmp[2504]*kernel[1]+tmp[2505]*kernel[2]+tmp[2603]*kernel[3]+tmp[2604]*kernel[4]+tmp[2605]*kernel[5]+tmp[2703]*kernel[6]+tmp[2704]*kernel[7]+tmp[2705]*kernel[8];
				ans[2605]<=tmp[2504]*kernel[0]+tmp[2505]*kernel[1]+tmp[2506]*kernel[2]+tmp[2604]*kernel[3]+tmp[2605]*kernel[4]+tmp[2606]*kernel[5]+tmp[2704]*kernel[6]+tmp[2705]*kernel[7]+tmp[2706]*kernel[8];
				ans[2606]<=tmp[2505]*kernel[0]+tmp[2506]*kernel[1]+tmp[2507]*kernel[2]+tmp[2605]*kernel[3]+tmp[2606]*kernel[4]+tmp[2607]*kernel[5]+tmp[2705]*kernel[6]+tmp[2706]*kernel[7]+tmp[2707]*kernel[8];
				ans[2607]<=tmp[2506]*kernel[0]+tmp[2507]*kernel[1]+tmp[2508]*kernel[2]+tmp[2606]*kernel[3]+tmp[2607]*kernel[4]+tmp[2608]*kernel[5]+tmp[2706]*kernel[6]+tmp[2707]*kernel[7]+tmp[2708]*kernel[8];
				ans[2608]<=tmp[2507]*kernel[0]+tmp[2508]*kernel[1]+tmp[2509]*kernel[2]+tmp[2607]*kernel[3]+tmp[2608]*kernel[4]+tmp[2609]*kernel[5]+tmp[2707]*kernel[6]+tmp[2708]*kernel[7]+tmp[2709]*kernel[8];
				ans[2609]<=tmp[2508]*kernel[0]+tmp[2509]*kernel[1]+tmp[2510]*kernel[2]+tmp[2608]*kernel[3]+tmp[2609]*kernel[4]+tmp[2610]*kernel[5]+tmp[2708]*kernel[6]+tmp[2709]*kernel[7]+tmp[2710]*kernel[8];
				ans[2610]<=tmp[2509]*kernel[0]+tmp[2510]*kernel[1]+tmp[2511]*kernel[2]+tmp[2609]*kernel[3]+tmp[2610]*kernel[4]+tmp[2611]*kernel[5]+tmp[2709]*kernel[6]+tmp[2710]*kernel[7]+tmp[2711]*kernel[8];
				ans[2611]<=tmp[2510]*kernel[0]+tmp[2511]*kernel[1]+tmp[2512]*kernel[2]+tmp[2610]*kernel[3]+tmp[2611]*kernel[4]+tmp[2612]*kernel[5]+tmp[2710]*kernel[6]+tmp[2711]*kernel[7]+tmp[2712]*kernel[8];
				ans[2612]<=tmp[2511]*kernel[0]+tmp[2512]*kernel[1]+tmp[2513]*kernel[2]+tmp[2611]*kernel[3]+tmp[2612]*kernel[4]+tmp[2613]*kernel[5]+tmp[2711]*kernel[6]+tmp[2712]*kernel[7]+tmp[2713]*kernel[8];
				ans[2613]<=tmp[2512]*kernel[0]+tmp[2513]*kernel[1]+tmp[2514]*kernel[2]+tmp[2612]*kernel[3]+tmp[2613]*kernel[4]+tmp[2614]*kernel[5]+tmp[2712]*kernel[6]+tmp[2713]*kernel[7]+tmp[2714]*kernel[8];
				ans[2614]<=tmp[2513]*kernel[0]+tmp[2514]*kernel[1]+tmp[2515]*kernel[2]+tmp[2613]*kernel[3]+tmp[2614]*kernel[4]+tmp[2615]*kernel[5]+tmp[2713]*kernel[6]+tmp[2714]*kernel[7]+tmp[2715]*kernel[8];
				ans[2615]<=tmp[2514]*kernel[0]+tmp[2515]*kernel[1]+tmp[2516]*kernel[2]+tmp[2614]*kernel[3]+tmp[2615]*kernel[4]+tmp[2616]*kernel[5]+tmp[2714]*kernel[6]+tmp[2715]*kernel[7]+tmp[2716]*kernel[8];
				ans[2616]<=tmp[2515]*kernel[0]+tmp[2516]*kernel[1]+tmp[2517]*kernel[2]+tmp[2615]*kernel[3]+tmp[2616]*kernel[4]+tmp[2617]*kernel[5]+tmp[2715]*kernel[6]+tmp[2716]*kernel[7]+tmp[2717]*kernel[8];
				ans[2617]<=tmp[2516]*kernel[0]+tmp[2517]*kernel[1]+tmp[2518]*kernel[2]+tmp[2616]*kernel[3]+tmp[2617]*kernel[4]+tmp[2618]*kernel[5]+tmp[2716]*kernel[6]+tmp[2717]*kernel[7]+tmp[2718]*kernel[8];
				ans[2618]<=tmp[2517]*kernel[0]+tmp[2518]*kernel[1]+tmp[2519]*kernel[2]+tmp[2617]*kernel[3]+tmp[2618]*kernel[4]+tmp[2619]*kernel[5]+tmp[2717]*kernel[6]+tmp[2718]*kernel[7]+tmp[2719]*kernel[8];
				ans[2619]<=tmp[2518]*kernel[0]+tmp[2519]*kernel[1]+tmp[2520]*kernel[2]+tmp[2618]*kernel[3]+tmp[2619]*kernel[4]+tmp[2620]*kernel[5]+tmp[2718]*kernel[6]+tmp[2719]*kernel[7]+tmp[2720]*kernel[8];
				ans[2620]<=tmp[2519]*kernel[0]+tmp[2520]*kernel[1]+tmp[2521]*kernel[2]+tmp[2619]*kernel[3]+tmp[2620]*kernel[4]+tmp[2621]*kernel[5]+tmp[2719]*kernel[6]+tmp[2720]*kernel[7]+tmp[2721]*kernel[8];
				ans[2621]<=tmp[2520]*kernel[0]+tmp[2521]*kernel[1]+tmp[2522]*kernel[2]+tmp[2620]*kernel[3]+tmp[2621]*kernel[4]+tmp[2622]*kernel[5]+tmp[2720]*kernel[6]+tmp[2721]*kernel[7]+tmp[2722]*kernel[8];
				ans[2622]<=tmp[2521]*kernel[0]+tmp[2522]*kernel[1]+tmp[2523]*kernel[2]+tmp[2621]*kernel[3]+tmp[2622]*kernel[4]+tmp[2623]*kernel[5]+tmp[2721]*kernel[6]+tmp[2722]*kernel[7]+tmp[2723]*kernel[8];
				ans[2623]<=tmp[2522]*kernel[0]+tmp[2523]*kernel[1]+tmp[2524]*kernel[2]+tmp[2622]*kernel[3]+tmp[2623]*kernel[4]+tmp[2624]*kernel[5]+tmp[2722]*kernel[6]+tmp[2723]*kernel[7]+tmp[2724]*kernel[8];
				ans[2624]<=tmp[2523]*kernel[0]+tmp[2524]*kernel[1]+tmp[2525]*kernel[2]+tmp[2623]*kernel[3]+tmp[2624]*kernel[4]+tmp[2625]*kernel[5]+tmp[2723]*kernel[6]+tmp[2724]*kernel[7]+tmp[2725]*kernel[8];
				ans[2625]<=tmp[2524]*kernel[0]+tmp[2525]*kernel[1]+tmp[2526]*kernel[2]+tmp[2624]*kernel[3]+tmp[2625]*kernel[4]+tmp[2626]*kernel[5]+tmp[2724]*kernel[6]+tmp[2725]*kernel[7]+tmp[2726]*kernel[8];
				ans[2626]<=tmp[2525]*kernel[0]+tmp[2526]*kernel[1]+tmp[2527]*kernel[2]+tmp[2625]*kernel[3]+tmp[2626]*kernel[4]+tmp[2627]*kernel[5]+tmp[2725]*kernel[6]+tmp[2726]*kernel[7]+tmp[2727]*kernel[8];
				ans[2627]<=tmp[2526]*kernel[0]+tmp[2527]*kernel[1]+tmp[2528]*kernel[2]+tmp[2626]*kernel[3]+tmp[2627]*kernel[4]+tmp[2628]*kernel[5]+tmp[2726]*kernel[6]+tmp[2727]*kernel[7]+tmp[2728]*kernel[8];
				ans[2628]<=tmp[2527]*kernel[0]+tmp[2528]*kernel[1]+tmp[2529]*kernel[2]+tmp[2627]*kernel[3]+tmp[2628]*kernel[4]+tmp[2629]*kernel[5]+tmp[2727]*kernel[6]+tmp[2728]*kernel[7]+tmp[2729]*kernel[8];
				ans[2629]<=tmp[2528]*kernel[0]+tmp[2529]*kernel[1]+tmp[2530]*kernel[2]+tmp[2628]*kernel[3]+tmp[2629]*kernel[4]+tmp[2630]*kernel[5]+tmp[2728]*kernel[6]+tmp[2729]*kernel[7]+tmp[2730]*kernel[8];
				ans[2630]<=tmp[2529]*kernel[0]+tmp[2530]*kernel[1]+tmp[2531]*kernel[2]+tmp[2629]*kernel[3]+tmp[2630]*kernel[4]+tmp[2631]*kernel[5]+tmp[2729]*kernel[6]+tmp[2730]*kernel[7]+tmp[2731]*kernel[8];
				ans[2631]<=tmp[2530]*kernel[0]+tmp[2531]*kernel[1]+tmp[2532]*kernel[2]+tmp[2630]*kernel[3]+tmp[2631]*kernel[4]+tmp[2632]*kernel[5]+tmp[2730]*kernel[6]+tmp[2731]*kernel[7]+tmp[2732]*kernel[8];
				ans[2632]<=tmp[2531]*kernel[0]+tmp[2532]*kernel[1]+tmp[2533]*kernel[2]+tmp[2631]*kernel[3]+tmp[2632]*kernel[4]+tmp[2633]*kernel[5]+tmp[2731]*kernel[6]+tmp[2732]*kernel[7]+tmp[2733]*kernel[8];
				ans[2633]<=tmp[2532]*kernel[0]+tmp[2533]*kernel[1]+tmp[2534]*kernel[2]+tmp[2632]*kernel[3]+tmp[2633]*kernel[4]+tmp[2634]*kernel[5]+tmp[2732]*kernel[6]+tmp[2733]*kernel[7]+tmp[2734]*kernel[8];
				ans[2634]<=tmp[2533]*kernel[0]+tmp[2534]*kernel[1]+tmp[2535]*kernel[2]+tmp[2633]*kernel[3]+tmp[2634]*kernel[4]+tmp[2635]*kernel[5]+tmp[2733]*kernel[6]+tmp[2734]*kernel[7]+tmp[2735]*kernel[8];
				ans[2635]<=tmp[2534]*kernel[0]+tmp[2535]*kernel[1]+tmp[2536]*kernel[2]+tmp[2634]*kernel[3]+tmp[2635]*kernel[4]+tmp[2636]*kernel[5]+tmp[2734]*kernel[6]+tmp[2735]*kernel[7]+tmp[2736]*kernel[8];
				ans[2636]<=tmp[2535]*kernel[0]+tmp[2536]*kernel[1]+tmp[2537]*kernel[2]+tmp[2635]*kernel[3]+tmp[2636]*kernel[4]+tmp[2637]*kernel[5]+tmp[2735]*kernel[6]+tmp[2736]*kernel[7]+tmp[2737]*kernel[8];
				ans[2637]<=tmp[2536]*kernel[0]+tmp[2537]*kernel[1]+tmp[2538]*kernel[2]+tmp[2636]*kernel[3]+tmp[2637]*kernel[4]+tmp[2638]*kernel[5]+tmp[2736]*kernel[6]+tmp[2737]*kernel[7]+tmp[2738]*kernel[8];
				ans[2638]<=tmp[2537]*kernel[0]+tmp[2538]*kernel[1]+tmp[2539]*kernel[2]+tmp[2637]*kernel[3]+tmp[2638]*kernel[4]+tmp[2639]*kernel[5]+tmp[2737]*kernel[6]+tmp[2738]*kernel[7]+tmp[2739]*kernel[8];
				ans[2639]<=tmp[2538]*kernel[0]+tmp[2539]*kernel[1]+tmp[2540]*kernel[2]+tmp[2638]*kernel[3]+tmp[2639]*kernel[4]+tmp[2640]*kernel[5]+tmp[2738]*kernel[6]+tmp[2739]*kernel[7]+tmp[2740]*kernel[8];
				ans[2640]<=tmp[2539]*kernel[0]+tmp[2540]*kernel[1]+tmp[2541]*kernel[2]+tmp[2639]*kernel[3]+tmp[2640]*kernel[4]+tmp[2641]*kernel[5]+tmp[2739]*kernel[6]+tmp[2740]*kernel[7]+tmp[2741]*kernel[8];
				ans[2641]<=tmp[2540]*kernel[0]+tmp[2541]*kernel[1]+tmp[2542]*kernel[2]+tmp[2640]*kernel[3]+tmp[2641]*kernel[4]+tmp[2642]*kernel[5]+tmp[2740]*kernel[6]+tmp[2741]*kernel[7]+tmp[2742]*kernel[8];
				ans[2642]<=tmp[2541]*kernel[0]+tmp[2542]*kernel[1]+tmp[2543]*kernel[2]+tmp[2641]*kernel[3]+tmp[2642]*kernel[4]+tmp[2643]*kernel[5]+tmp[2741]*kernel[6]+tmp[2742]*kernel[7]+tmp[2743]*kernel[8];
				ans[2643]<=tmp[2542]*kernel[0]+tmp[2543]*kernel[1]+tmp[2544]*kernel[2]+tmp[2642]*kernel[3]+tmp[2643]*kernel[4]+tmp[2644]*kernel[5]+tmp[2742]*kernel[6]+tmp[2743]*kernel[7]+tmp[2744]*kernel[8];
				ans[2644]<=tmp[2543]*kernel[0]+tmp[2544]*kernel[1]+tmp[2545]*kernel[2]+tmp[2643]*kernel[3]+tmp[2644]*kernel[4]+tmp[2645]*kernel[5]+tmp[2743]*kernel[6]+tmp[2744]*kernel[7]+tmp[2745]*kernel[8];
				ans[2645]<=tmp[2544]*kernel[0]+tmp[2545]*kernel[1]+tmp[2546]*kernel[2]+tmp[2644]*kernel[3]+tmp[2645]*kernel[4]+tmp[2646]*kernel[5]+tmp[2744]*kernel[6]+tmp[2745]*kernel[7]+tmp[2746]*kernel[8];
				ans[2646]<=tmp[2545]*kernel[0]+tmp[2546]*kernel[1]+tmp[2547]*kernel[2]+tmp[2645]*kernel[3]+tmp[2646]*kernel[4]+tmp[2647]*kernel[5]+tmp[2745]*kernel[6]+tmp[2746]*kernel[7]+tmp[2747]*kernel[8];
				ans[2647]<=tmp[2546]*kernel[0]+tmp[2547]*kernel[1]+tmp[2548]*kernel[2]+tmp[2646]*kernel[3]+tmp[2647]*kernel[4]+tmp[2648]*kernel[5]+tmp[2746]*kernel[6]+tmp[2747]*kernel[7]+tmp[2748]*kernel[8];
				ans[2648]<=tmp[2547]*kernel[0]+tmp[2548]*kernel[1]+tmp[2549]*kernel[2]+tmp[2647]*kernel[3]+tmp[2648]*kernel[4]+tmp[2649]*kernel[5]+tmp[2747]*kernel[6]+tmp[2748]*kernel[7]+tmp[2749]*kernel[8];
				ans[2649]<=tmp[2548]*kernel[0]+tmp[2549]*kernel[1]+tmp[2550]*kernel[2]+tmp[2648]*kernel[3]+tmp[2649]*kernel[4]+tmp[2650]*kernel[5]+tmp[2748]*kernel[6]+tmp[2749]*kernel[7]+tmp[2750]*kernel[8];
				ans[2650]<=tmp[2549]*kernel[0]+tmp[2550]*kernel[1]+tmp[2551]*kernel[2]+tmp[2649]*kernel[3]+tmp[2650]*kernel[4]+tmp[2651]*kernel[5]+tmp[2749]*kernel[6]+tmp[2750]*kernel[7]+tmp[2751]*kernel[8];
				ans[2651]<=tmp[2550]*kernel[0]+tmp[2551]*kernel[1]+tmp[2552]*kernel[2]+tmp[2650]*kernel[3]+tmp[2651]*kernel[4]+tmp[2652]*kernel[5]+tmp[2750]*kernel[6]+tmp[2751]*kernel[7]+tmp[2752]*kernel[8];
				ans[2652]<=tmp[2551]*kernel[0]+tmp[2552]*kernel[1]+tmp[2553]*kernel[2]+tmp[2651]*kernel[3]+tmp[2652]*kernel[4]+tmp[2653]*kernel[5]+tmp[2751]*kernel[6]+tmp[2752]*kernel[7]+tmp[2753]*kernel[8];
				ans[2653]<=tmp[2552]*kernel[0]+tmp[2553]*kernel[1]+tmp[2554]*kernel[2]+tmp[2652]*kernel[3]+tmp[2653]*kernel[4]+tmp[2654]*kernel[5]+tmp[2752]*kernel[6]+tmp[2753]*kernel[7]+tmp[2754]*kernel[8];
				ans[2654]<=tmp[2553]*kernel[0]+tmp[2554]*kernel[1]+tmp[2555]*kernel[2]+tmp[2653]*kernel[3]+tmp[2654]*kernel[4]+tmp[2655]*kernel[5]+tmp[2753]*kernel[6]+tmp[2754]*kernel[7]+tmp[2755]*kernel[8];
				ans[2655]<=tmp[2554]*kernel[0]+tmp[2555]*kernel[1]+tmp[2556]*kernel[2]+tmp[2654]*kernel[3]+tmp[2655]*kernel[4]+tmp[2656]*kernel[5]+tmp[2754]*kernel[6]+tmp[2755]*kernel[7]+tmp[2756]*kernel[8];
				ans[2656]<=tmp[2555]*kernel[0]+tmp[2556]*kernel[1]+tmp[2557]*kernel[2]+tmp[2655]*kernel[3]+tmp[2656]*kernel[4]+tmp[2657]*kernel[5]+tmp[2755]*kernel[6]+tmp[2756]*kernel[7]+tmp[2757]*kernel[8];
				ans[2657]<=tmp[2556]*kernel[0]+tmp[2557]*kernel[1]+tmp[2558]*kernel[2]+tmp[2656]*kernel[3]+tmp[2657]*kernel[4]+tmp[2658]*kernel[5]+tmp[2756]*kernel[6]+tmp[2757]*kernel[7]+tmp[2758]*kernel[8];
				ans[2658]<=tmp[2557]*kernel[0]+tmp[2558]*kernel[1]+tmp[2559]*kernel[2]+tmp[2657]*kernel[3]+tmp[2658]*kernel[4]+tmp[2659]*kernel[5]+tmp[2757]*kernel[6]+tmp[2758]*kernel[7]+tmp[2759]*kernel[8];
				ans[2659]<=tmp[2558]*kernel[0]+tmp[2559]*kernel[1]+tmp[2560]*kernel[2]+tmp[2658]*kernel[3]+tmp[2659]*kernel[4]+tmp[2660]*kernel[5]+tmp[2758]*kernel[6]+tmp[2759]*kernel[7]+tmp[2760]*kernel[8];
				ans[2660]<=tmp[2559]*kernel[0]+tmp[2560]*kernel[1]+tmp[2561]*kernel[2]+tmp[2659]*kernel[3]+tmp[2660]*kernel[4]+tmp[2661]*kernel[5]+tmp[2759]*kernel[6]+tmp[2760]*kernel[7]+tmp[2761]*kernel[8];
				ans[2661]<=tmp[2560]*kernel[0]+tmp[2561]*kernel[1]+tmp[2562]*kernel[2]+tmp[2660]*kernel[3]+tmp[2661]*kernel[4]+tmp[2662]*kernel[5]+tmp[2760]*kernel[6]+tmp[2761]*kernel[7]+tmp[2762]*kernel[8];
				ans[2662]<=tmp[2561]*kernel[0]+tmp[2562]*kernel[1]+tmp[2563]*kernel[2]+tmp[2661]*kernel[3]+tmp[2662]*kernel[4]+tmp[2663]*kernel[5]+tmp[2761]*kernel[6]+tmp[2762]*kernel[7]+tmp[2763]*kernel[8];
				ans[2663]<=tmp[2562]*kernel[0]+tmp[2563]*kernel[1]+tmp[2564]*kernel[2]+tmp[2662]*kernel[3]+tmp[2663]*kernel[4]+tmp[2664]*kernel[5]+tmp[2762]*kernel[6]+tmp[2763]*kernel[7]+tmp[2764]*kernel[8];
				ans[2664]<=tmp[2563]*kernel[0]+tmp[2564]*kernel[1]+tmp[2565]*kernel[2]+tmp[2663]*kernel[3]+tmp[2664]*kernel[4]+tmp[2665]*kernel[5]+tmp[2763]*kernel[6]+tmp[2764]*kernel[7]+tmp[2765]*kernel[8];
				ans[2665]<=tmp[2564]*kernel[0]+tmp[2565]*kernel[1]+tmp[2566]*kernel[2]+tmp[2664]*kernel[3]+tmp[2665]*kernel[4]+tmp[2666]*kernel[5]+tmp[2764]*kernel[6]+tmp[2765]*kernel[7]+tmp[2766]*kernel[8];
				ans[2666]<=tmp[2565]*kernel[0]+tmp[2566]*kernel[1]+tmp[2567]*kernel[2]+tmp[2665]*kernel[3]+tmp[2666]*kernel[4]+tmp[2667]*kernel[5]+tmp[2765]*kernel[6]+tmp[2766]*kernel[7]+tmp[2767]*kernel[8];
				ans[2667]<=tmp[2566]*kernel[0]+tmp[2567]*kernel[1]+tmp[2568]*kernel[2]+tmp[2666]*kernel[3]+tmp[2667]*kernel[4]+tmp[2668]*kernel[5]+tmp[2766]*kernel[6]+tmp[2767]*kernel[7]+tmp[2768]*kernel[8];
				ans[2668]<=tmp[2567]*kernel[0]+tmp[2568]*kernel[1]+tmp[2569]*kernel[2]+tmp[2667]*kernel[3]+tmp[2668]*kernel[4]+tmp[2669]*kernel[5]+tmp[2767]*kernel[6]+tmp[2768]*kernel[7]+tmp[2769]*kernel[8];
				ans[2669]<=tmp[2568]*kernel[0]+tmp[2569]*kernel[1]+tmp[2570]*kernel[2]+tmp[2668]*kernel[3]+tmp[2669]*kernel[4]+tmp[2670]*kernel[5]+tmp[2768]*kernel[6]+tmp[2769]*kernel[7]+tmp[2770]*kernel[8];
				ans[2670]<=tmp[2569]*kernel[0]+tmp[2570]*kernel[1]+tmp[2571]*kernel[2]+tmp[2669]*kernel[3]+tmp[2670]*kernel[4]+tmp[2671]*kernel[5]+tmp[2769]*kernel[6]+tmp[2770]*kernel[7]+tmp[2771]*kernel[8];
				ans[2671]<=tmp[2570]*kernel[0]+tmp[2571]*kernel[1]+tmp[2572]*kernel[2]+tmp[2670]*kernel[3]+tmp[2671]*kernel[4]+tmp[2672]*kernel[5]+tmp[2770]*kernel[6]+tmp[2771]*kernel[7]+tmp[2772]*kernel[8];
				ans[2672]<=tmp[2571]*kernel[0]+tmp[2572]*kernel[1]+tmp[2573]*kernel[2]+tmp[2671]*kernel[3]+tmp[2672]*kernel[4]+tmp[2673]*kernel[5]+tmp[2771]*kernel[6]+tmp[2772]*kernel[7]+tmp[2773]*kernel[8];
				ans[2673]<=tmp[2572]*kernel[0]+tmp[2573]*kernel[1]+tmp[2574]*kernel[2]+tmp[2672]*kernel[3]+tmp[2673]*kernel[4]+tmp[2674]*kernel[5]+tmp[2772]*kernel[6]+tmp[2773]*kernel[7]+tmp[2774]*kernel[8];
				ans[2674]<=tmp[2573]*kernel[0]+tmp[2574]*kernel[1]+tmp[2575]*kernel[2]+tmp[2673]*kernel[3]+tmp[2674]*kernel[4]+tmp[2675]*kernel[5]+tmp[2773]*kernel[6]+tmp[2774]*kernel[7]+tmp[2775]*kernel[8];
				ans[2675]<=tmp[2574]*kernel[0]+tmp[2575]*kernel[1]+tmp[2576]*kernel[2]+tmp[2674]*kernel[3]+tmp[2675]*kernel[4]+tmp[2676]*kernel[5]+tmp[2774]*kernel[6]+tmp[2775]*kernel[7]+tmp[2776]*kernel[8];
				ans[2676]<=tmp[2575]*kernel[0]+tmp[2576]*kernel[1]+tmp[2577]*kernel[2]+tmp[2675]*kernel[3]+tmp[2676]*kernel[4]+tmp[2677]*kernel[5]+tmp[2775]*kernel[6]+tmp[2776]*kernel[7]+tmp[2777]*kernel[8];
				ans[2677]<=tmp[2576]*kernel[0]+tmp[2577]*kernel[1]+tmp[2578]*kernel[2]+tmp[2676]*kernel[3]+tmp[2677]*kernel[4]+tmp[2678]*kernel[5]+tmp[2776]*kernel[6]+tmp[2777]*kernel[7]+tmp[2778]*kernel[8];
				ans[2678]<=tmp[2577]*kernel[0]+tmp[2578]*kernel[1]+tmp[2579]*kernel[2]+tmp[2677]*kernel[3]+tmp[2678]*kernel[4]+tmp[2679]*kernel[5]+tmp[2777]*kernel[6]+tmp[2778]*kernel[7]+tmp[2779]*kernel[8];
				ans[2679]<=tmp[2578]*kernel[0]+tmp[2579]*kernel[1]+tmp[2580]*kernel[2]+tmp[2678]*kernel[3]+tmp[2679]*kernel[4]+tmp[2680]*kernel[5]+tmp[2778]*kernel[6]+tmp[2779]*kernel[7]+tmp[2780]*kernel[8];
				ans[2680]<=tmp[2579]*kernel[0]+tmp[2580]*kernel[1]+tmp[2581]*kernel[2]+tmp[2679]*kernel[3]+tmp[2680]*kernel[4]+tmp[2681]*kernel[5]+tmp[2779]*kernel[6]+tmp[2780]*kernel[7]+tmp[2781]*kernel[8];
				ans[2681]<=tmp[2580]*kernel[0]+tmp[2581]*kernel[1]+tmp[2582]*kernel[2]+tmp[2680]*kernel[3]+tmp[2681]*kernel[4]+tmp[2682]*kernel[5]+tmp[2780]*kernel[6]+tmp[2781]*kernel[7]+tmp[2782]*kernel[8];
				ans[2682]<=tmp[2581]*kernel[0]+tmp[2582]*kernel[1]+tmp[2583]*kernel[2]+tmp[2681]*kernel[3]+tmp[2682]*kernel[4]+tmp[2683]*kernel[5]+tmp[2781]*kernel[6]+tmp[2782]*kernel[7]+tmp[2783]*kernel[8];
				ans[2683]<=tmp[2582]*kernel[0]+tmp[2583]*kernel[1]+tmp[2584]*kernel[2]+tmp[2682]*kernel[3]+tmp[2683]*kernel[4]+tmp[2684]*kernel[5]+tmp[2782]*kernel[6]+tmp[2783]*kernel[7]+tmp[2784]*kernel[8];
				ans[2684]<=tmp[2583]*kernel[0]+tmp[2584]*kernel[1]+tmp[2585]*kernel[2]+tmp[2683]*kernel[3]+tmp[2684]*kernel[4]+tmp[2685]*kernel[5]+tmp[2783]*kernel[6]+tmp[2784]*kernel[7]+tmp[2785]*kernel[8];
				ans[2685]<=tmp[2584]*kernel[0]+tmp[2585]*kernel[1]+tmp[2586]*kernel[2]+tmp[2684]*kernel[3]+tmp[2685]*kernel[4]+tmp[2686]*kernel[5]+tmp[2784]*kernel[6]+tmp[2785]*kernel[7]+tmp[2786]*kernel[8];
				ans[2686]<=tmp[2585]*kernel[0]+tmp[2586]*kernel[1]+tmp[2587]*kernel[2]+tmp[2685]*kernel[3]+tmp[2686]*kernel[4]+tmp[2687]*kernel[5]+tmp[2785]*kernel[6]+tmp[2786]*kernel[7]+tmp[2787]*kernel[8];
				ans[2687]<=tmp[2586]*kernel[0]+tmp[2587]*kernel[1]+tmp[2588]*kernel[2]+tmp[2686]*kernel[3]+tmp[2687]*kernel[4]+tmp[2688]*kernel[5]+tmp[2786]*kernel[6]+tmp[2787]*kernel[7]+tmp[2788]*kernel[8];
				ans[2688]<=tmp[2587]*kernel[0]+tmp[2588]*kernel[1]+tmp[2589]*kernel[2]+tmp[2687]*kernel[3]+tmp[2688]*kernel[4]+tmp[2689]*kernel[5]+tmp[2787]*kernel[6]+tmp[2788]*kernel[7]+tmp[2789]*kernel[8];
				ans[2689]<=tmp[2588]*kernel[0]+tmp[2589]*kernel[1]+tmp[2590]*kernel[2]+tmp[2688]*kernel[3]+tmp[2689]*kernel[4]+tmp[2690]*kernel[5]+tmp[2788]*kernel[6]+tmp[2789]*kernel[7]+tmp[2790]*kernel[8];
				ans[2690]<=tmp[2589]*kernel[0]+tmp[2590]*kernel[1]+tmp[2591]*kernel[2]+tmp[2689]*kernel[3]+tmp[2690]*kernel[4]+tmp[2691]*kernel[5]+tmp[2789]*kernel[6]+tmp[2790]*kernel[7]+tmp[2791]*kernel[8];
				ans[2691]<=tmp[2590]*kernel[0]+tmp[2591]*kernel[1]+tmp[2592]*kernel[2]+tmp[2690]*kernel[3]+tmp[2691]*kernel[4]+tmp[2692]*kernel[5]+tmp[2790]*kernel[6]+tmp[2791]*kernel[7]+tmp[2792]*kernel[8];
				ans[2692]<=tmp[2591]*kernel[0]+tmp[2592]*kernel[1]+tmp[2593]*kernel[2]+tmp[2691]*kernel[3]+tmp[2692]*kernel[4]+tmp[2693]*kernel[5]+tmp[2791]*kernel[6]+tmp[2792]*kernel[7]+tmp[2793]*kernel[8];
				ans[2693]<=tmp[2592]*kernel[0]+tmp[2593]*kernel[1]+tmp[2594]*kernel[2]+tmp[2692]*kernel[3]+tmp[2693]*kernel[4]+tmp[2694]*kernel[5]+tmp[2792]*kernel[6]+tmp[2793]*kernel[7]+tmp[2794]*kernel[8];
				ans[2694]<=tmp[2593]*kernel[0]+tmp[2594]*kernel[1]+tmp[2595]*kernel[2]+tmp[2693]*kernel[3]+tmp[2694]*kernel[4]+tmp[2695]*kernel[5]+tmp[2793]*kernel[6]+tmp[2794]*kernel[7]+tmp[2795]*kernel[8];
				ans[2695]<=tmp[2594]*kernel[0]+tmp[2595]*kernel[1]+tmp[2596]*kernel[2]+tmp[2694]*kernel[3]+tmp[2695]*kernel[4]+tmp[2696]*kernel[5]+tmp[2794]*kernel[6]+tmp[2795]*kernel[7]+tmp[2796]*kernel[8];
				ans[2696]<=tmp[2595]*kernel[0]+tmp[2596]*kernel[1]+tmp[2597]*kernel[2]+tmp[2695]*kernel[3]+tmp[2696]*kernel[4]+tmp[2697]*kernel[5]+tmp[2795]*kernel[6]+tmp[2796]*kernel[7]+tmp[2797]*kernel[8];
				ans[2697]<=tmp[2596]*kernel[0]+tmp[2597]*kernel[1]+tmp[2598]*kernel[2]+tmp[2696]*kernel[3]+tmp[2697]*kernel[4]+tmp[2698]*kernel[5]+tmp[2796]*kernel[6]+tmp[2797]*kernel[7]+tmp[2798]*kernel[8];
				ans[2698]<=tmp[2597]*kernel[0]+tmp[2598]*kernel[1]+tmp[2599]*kernel[2]+tmp[2697]*kernel[3]+tmp[2698]*kernel[4]+tmp[2699]*kernel[5]+tmp[2797]*kernel[6]+tmp[2798]*kernel[7]+tmp[2799]*kernel[8];
				ans[2699]<=tmp[2598]*kernel[0]+tmp[2599]*kernel[1]+tmp[2698]*kernel[3]+tmp[2699]*kernel[4]+tmp[2798]*kernel[6]+tmp[2799]*kernel[7];
				ans[2700]<=tmp[2600]*kernel[1]+tmp[2601]*kernel[2]+tmp[2700]*kernel[4]+tmp[2701]*kernel[5]+tmp[2800]*kernel[7]+tmp[2801]*kernel[8];
				ans[2701]<=tmp[2600]*kernel[0]+tmp[2601]*kernel[1]+tmp[2602]*kernel[2]+tmp[2700]*kernel[3]+tmp[2701]*kernel[4]+tmp[2702]*kernel[5]+tmp[2800]*kernel[6]+tmp[2801]*kernel[7]+tmp[2802]*kernel[8];
				ans[2702]<=tmp[2601]*kernel[0]+tmp[2602]*kernel[1]+tmp[2603]*kernel[2]+tmp[2701]*kernel[3]+tmp[2702]*kernel[4]+tmp[2703]*kernel[5]+tmp[2801]*kernel[6]+tmp[2802]*kernel[7]+tmp[2803]*kernel[8];
				ans[2703]<=tmp[2602]*kernel[0]+tmp[2603]*kernel[1]+tmp[2604]*kernel[2]+tmp[2702]*kernel[3]+tmp[2703]*kernel[4]+tmp[2704]*kernel[5]+tmp[2802]*kernel[6]+tmp[2803]*kernel[7]+tmp[2804]*kernel[8];
				ans[2704]<=tmp[2603]*kernel[0]+tmp[2604]*kernel[1]+tmp[2605]*kernel[2]+tmp[2703]*kernel[3]+tmp[2704]*kernel[4]+tmp[2705]*kernel[5]+tmp[2803]*kernel[6]+tmp[2804]*kernel[7]+tmp[2805]*kernel[8];
				ans[2705]<=tmp[2604]*kernel[0]+tmp[2605]*kernel[1]+tmp[2606]*kernel[2]+tmp[2704]*kernel[3]+tmp[2705]*kernel[4]+tmp[2706]*kernel[5]+tmp[2804]*kernel[6]+tmp[2805]*kernel[7]+tmp[2806]*kernel[8];
				ans[2706]<=tmp[2605]*kernel[0]+tmp[2606]*kernel[1]+tmp[2607]*kernel[2]+tmp[2705]*kernel[3]+tmp[2706]*kernel[4]+tmp[2707]*kernel[5]+tmp[2805]*kernel[6]+tmp[2806]*kernel[7]+tmp[2807]*kernel[8];
				ans[2707]<=tmp[2606]*kernel[0]+tmp[2607]*kernel[1]+tmp[2608]*kernel[2]+tmp[2706]*kernel[3]+tmp[2707]*kernel[4]+tmp[2708]*kernel[5]+tmp[2806]*kernel[6]+tmp[2807]*kernel[7]+tmp[2808]*kernel[8];
				ans[2708]<=tmp[2607]*kernel[0]+tmp[2608]*kernel[1]+tmp[2609]*kernel[2]+tmp[2707]*kernel[3]+tmp[2708]*kernel[4]+tmp[2709]*kernel[5]+tmp[2807]*kernel[6]+tmp[2808]*kernel[7]+tmp[2809]*kernel[8];
				ans[2709]<=tmp[2608]*kernel[0]+tmp[2609]*kernel[1]+tmp[2610]*kernel[2]+tmp[2708]*kernel[3]+tmp[2709]*kernel[4]+tmp[2710]*kernel[5]+tmp[2808]*kernel[6]+tmp[2809]*kernel[7]+tmp[2810]*kernel[8];
				ans[2710]<=tmp[2609]*kernel[0]+tmp[2610]*kernel[1]+tmp[2611]*kernel[2]+tmp[2709]*kernel[3]+tmp[2710]*kernel[4]+tmp[2711]*kernel[5]+tmp[2809]*kernel[6]+tmp[2810]*kernel[7]+tmp[2811]*kernel[8];
				ans[2711]<=tmp[2610]*kernel[0]+tmp[2611]*kernel[1]+tmp[2612]*kernel[2]+tmp[2710]*kernel[3]+tmp[2711]*kernel[4]+tmp[2712]*kernel[5]+tmp[2810]*kernel[6]+tmp[2811]*kernel[7]+tmp[2812]*kernel[8];
				ans[2712]<=tmp[2611]*kernel[0]+tmp[2612]*kernel[1]+tmp[2613]*kernel[2]+tmp[2711]*kernel[3]+tmp[2712]*kernel[4]+tmp[2713]*kernel[5]+tmp[2811]*kernel[6]+tmp[2812]*kernel[7]+tmp[2813]*kernel[8];
				ans[2713]<=tmp[2612]*kernel[0]+tmp[2613]*kernel[1]+tmp[2614]*kernel[2]+tmp[2712]*kernel[3]+tmp[2713]*kernel[4]+tmp[2714]*kernel[5]+tmp[2812]*kernel[6]+tmp[2813]*kernel[7]+tmp[2814]*kernel[8];
				ans[2714]<=tmp[2613]*kernel[0]+tmp[2614]*kernel[1]+tmp[2615]*kernel[2]+tmp[2713]*kernel[3]+tmp[2714]*kernel[4]+tmp[2715]*kernel[5]+tmp[2813]*kernel[6]+tmp[2814]*kernel[7]+tmp[2815]*kernel[8];
				ans[2715]<=tmp[2614]*kernel[0]+tmp[2615]*kernel[1]+tmp[2616]*kernel[2]+tmp[2714]*kernel[3]+tmp[2715]*kernel[4]+tmp[2716]*kernel[5]+tmp[2814]*kernel[6]+tmp[2815]*kernel[7]+tmp[2816]*kernel[8];
				ans[2716]<=tmp[2615]*kernel[0]+tmp[2616]*kernel[1]+tmp[2617]*kernel[2]+tmp[2715]*kernel[3]+tmp[2716]*kernel[4]+tmp[2717]*kernel[5]+tmp[2815]*kernel[6]+tmp[2816]*kernel[7]+tmp[2817]*kernel[8];
				ans[2717]<=tmp[2616]*kernel[0]+tmp[2617]*kernel[1]+tmp[2618]*kernel[2]+tmp[2716]*kernel[3]+tmp[2717]*kernel[4]+tmp[2718]*kernel[5]+tmp[2816]*kernel[6]+tmp[2817]*kernel[7]+tmp[2818]*kernel[8];
				ans[2718]<=tmp[2617]*kernel[0]+tmp[2618]*kernel[1]+tmp[2619]*kernel[2]+tmp[2717]*kernel[3]+tmp[2718]*kernel[4]+tmp[2719]*kernel[5]+tmp[2817]*kernel[6]+tmp[2818]*kernel[7]+tmp[2819]*kernel[8];
				ans[2719]<=tmp[2618]*kernel[0]+tmp[2619]*kernel[1]+tmp[2620]*kernel[2]+tmp[2718]*kernel[3]+tmp[2719]*kernel[4]+tmp[2720]*kernel[5]+tmp[2818]*kernel[6]+tmp[2819]*kernel[7]+tmp[2820]*kernel[8];
				ans[2720]<=tmp[2619]*kernel[0]+tmp[2620]*kernel[1]+tmp[2621]*kernel[2]+tmp[2719]*kernel[3]+tmp[2720]*kernel[4]+tmp[2721]*kernel[5]+tmp[2819]*kernel[6]+tmp[2820]*kernel[7]+tmp[2821]*kernel[8];
				ans[2721]<=tmp[2620]*kernel[0]+tmp[2621]*kernel[1]+tmp[2622]*kernel[2]+tmp[2720]*kernel[3]+tmp[2721]*kernel[4]+tmp[2722]*kernel[5]+tmp[2820]*kernel[6]+tmp[2821]*kernel[7]+tmp[2822]*kernel[8];
				ans[2722]<=tmp[2621]*kernel[0]+tmp[2622]*kernel[1]+tmp[2623]*kernel[2]+tmp[2721]*kernel[3]+tmp[2722]*kernel[4]+tmp[2723]*kernel[5]+tmp[2821]*kernel[6]+tmp[2822]*kernel[7]+tmp[2823]*kernel[8];
				ans[2723]<=tmp[2622]*kernel[0]+tmp[2623]*kernel[1]+tmp[2624]*kernel[2]+tmp[2722]*kernel[3]+tmp[2723]*kernel[4]+tmp[2724]*kernel[5]+tmp[2822]*kernel[6]+tmp[2823]*kernel[7]+tmp[2824]*kernel[8];
				ans[2724]<=tmp[2623]*kernel[0]+tmp[2624]*kernel[1]+tmp[2625]*kernel[2]+tmp[2723]*kernel[3]+tmp[2724]*kernel[4]+tmp[2725]*kernel[5]+tmp[2823]*kernel[6]+tmp[2824]*kernel[7]+tmp[2825]*kernel[8];
				ans[2725]<=tmp[2624]*kernel[0]+tmp[2625]*kernel[1]+tmp[2626]*kernel[2]+tmp[2724]*kernel[3]+tmp[2725]*kernel[4]+tmp[2726]*kernel[5]+tmp[2824]*kernel[6]+tmp[2825]*kernel[7]+tmp[2826]*kernel[8];
				ans[2726]<=tmp[2625]*kernel[0]+tmp[2626]*kernel[1]+tmp[2627]*kernel[2]+tmp[2725]*kernel[3]+tmp[2726]*kernel[4]+tmp[2727]*kernel[5]+tmp[2825]*kernel[6]+tmp[2826]*kernel[7]+tmp[2827]*kernel[8];
				ans[2727]<=tmp[2626]*kernel[0]+tmp[2627]*kernel[1]+tmp[2628]*kernel[2]+tmp[2726]*kernel[3]+tmp[2727]*kernel[4]+tmp[2728]*kernel[5]+tmp[2826]*kernel[6]+tmp[2827]*kernel[7]+tmp[2828]*kernel[8];
				ans[2728]<=tmp[2627]*kernel[0]+tmp[2628]*kernel[1]+tmp[2629]*kernel[2]+tmp[2727]*kernel[3]+tmp[2728]*kernel[4]+tmp[2729]*kernel[5]+tmp[2827]*kernel[6]+tmp[2828]*kernel[7]+tmp[2829]*kernel[8];
				ans[2729]<=tmp[2628]*kernel[0]+tmp[2629]*kernel[1]+tmp[2630]*kernel[2]+tmp[2728]*kernel[3]+tmp[2729]*kernel[4]+tmp[2730]*kernel[5]+tmp[2828]*kernel[6]+tmp[2829]*kernel[7]+tmp[2830]*kernel[8];
				ans[2730]<=tmp[2629]*kernel[0]+tmp[2630]*kernel[1]+tmp[2631]*kernel[2]+tmp[2729]*kernel[3]+tmp[2730]*kernel[4]+tmp[2731]*kernel[5]+tmp[2829]*kernel[6]+tmp[2830]*kernel[7]+tmp[2831]*kernel[8];
				ans[2731]<=tmp[2630]*kernel[0]+tmp[2631]*kernel[1]+tmp[2632]*kernel[2]+tmp[2730]*kernel[3]+tmp[2731]*kernel[4]+tmp[2732]*kernel[5]+tmp[2830]*kernel[6]+tmp[2831]*kernel[7]+tmp[2832]*kernel[8];
				ans[2732]<=tmp[2631]*kernel[0]+tmp[2632]*kernel[1]+tmp[2633]*kernel[2]+tmp[2731]*kernel[3]+tmp[2732]*kernel[4]+tmp[2733]*kernel[5]+tmp[2831]*kernel[6]+tmp[2832]*kernel[7]+tmp[2833]*kernel[8];
				ans[2733]<=tmp[2632]*kernel[0]+tmp[2633]*kernel[1]+tmp[2634]*kernel[2]+tmp[2732]*kernel[3]+tmp[2733]*kernel[4]+tmp[2734]*kernel[5]+tmp[2832]*kernel[6]+tmp[2833]*kernel[7]+tmp[2834]*kernel[8];
				ans[2734]<=tmp[2633]*kernel[0]+tmp[2634]*kernel[1]+tmp[2635]*kernel[2]+tmp[2733]*kernel[3]+tmp[2734]*kernel[4]+tmp[2735]*kernel[5]+tmp[2833]*kernel[6]+tmp[2834]*kernel[7]+tmp[2835]*kernel[8];
				ans[2735]<=tmp[2634]*kernel[0]+tmp[2635]*kernel[1]+tmp[2636]*kernel[2]+tmp[2734]*kernel[3]+tmp[2735]*kernel[4]+tmp[2736]*kernel[5]+tmp[2834]*kernel[6]+tmp[2835]*kernel[7]+tmp[2836]*kernel[8];
				ans[2736]<=tmp[2635]*kernel[0]+tmp[2636]*kernel[1]+tmp[2637]*kernel[2]+tmp[2735]*kernel[3]+tmp[2736]*kernel[4]+tmp[2737]*kernel[5]+tmp[2835]*kernel[6]+tmp[2836]*kernel[7]+tmp[2837]*kernel[8];
				ans[2737]<=tmp[2636]*kernel[0]+tmp[2637]*kernel[1]+tmp[2638]*kernel[2]+tmp[2736]*kernel[3]+tmp[2737]*kernel[4]+tmp[2738]*kernel[5]+tmp[2836]*kernel[6]+tmp[2837]*kernel[7]+tmp[2838]*kernel[8];
				ans[2738]<=tmp[2637]*kernel[0]+tmp[2638]*kernel[1]+tmp[2639]*kernel[2]+tmp[2737]*kernel[3]+tmp[2738]*kernel[4]+tmp[2739]*kernel[5]+tmp[2837]*kernel[6]+tmp[2838]*kernel[7]+tmp[2839]*kernel[8];
				ans[2739]<=tmp[2638]*kernel[0]+tmp[2639]*kernel[1]+tmp[2640]*kernel[2]+tmp[2738]*kernel[3]+tmp[2739]*kernel[4]+tmp[2740]*kernel[5]+tmp[2838]*kernel[6]+tmp[2839]*kernel[7]+tmp[2840]*kernel[8];
				ans[2740]<=tmp[2639]*kernel[0]+tmp[2640]*kernel[1]+tmp[2641]*kernel[2]+tmp[2739]*kernel[3]+tmp[2740]*kernel[4]+tmp[2741]*kernel[5]+tmp[2839]*kernel[6]+tmp[2840]*kernel[7]+tmp[2841]*kernel[8];
				ans[2741]<=tmp[2640]*kernel[0]+tmp[2641]*kernel[1]+tmp[2642]*kernel[2]+tmp[2740]*kernel[3]+tmp[2741]*kernel[4]+tmp[2742]*kernel[5]+tmp[2840]*kernel[6]+tmp[2841]*kernel[7]+tmp[2842]*kernel[8];
				ans[2742]<=tmp[2641]*kernel[0]+tmp[2642]*kernel[1]+tmp[2643]*kernel[2]+tmp[2741]*kernel[3]+tmp[2742]*kernel[4]+tmp[2743]*kernel[5]+tmp[2841]*kernel[6]+tmp[2842]*kernel[7]+tmp[2843]*kernel[8];
				ans[2743]<=tmp[2642]*kernel[0]+tmp[2643]*kernel[1]+tmp[2644]*kernel[2]+tmp[2742]*kernel[3]+tmp[2743]*kernel[4]+tmp[2744]*kernel[5]+tmp[2842]*kernel[6]+tmp[2843]*kernel[7]+tmp[2844]*kernel[8];
				ans[2744]<=tmp[2643]*kernel[0]+tmp[2644]*kernel[1]+tmp[2645]*kernel[2]+tmp[2743]*kernel[3]+tmp[2744]*kernel[4]+tmp[2745]*kernel[5]+tmp[2843]*kernel[6]+tmp[2844]*kernel[7]+tmp[2845]*kernel[8];
				ans[2745]<=tmp[2644]*kernel[0]+tmp[2645]*kernel[1]+tmp[2646]*kernel[2]+tmp[2744]*kernel[3]+tmp[2745]*kernel[4]+tmp[2746]*kernel[5]+tmp[2844]*kernel[6]+tmp[2845]*kernel[7]+tmp[2846]*kernel[8];
				ans[2746]<=tmp[2645]*kernel[0]+tmp[2646]*kernel[1]+tmp[2647]*kernel[2]+tmp[2745]*kernel[3]+tmp[2746]*kernel[4]+tmp[2747]*kernel[5]+tmp[2845]*kernel[6]+tmp[2846]*kernel[7]+tmp[2847]*kernel[8];
				ans[2747]<=tmp[2646]*kernel[0]+tmp[2647]*kernel[1]+tmp[2648]*kernel[2]+tmp[2746]*kernel[3]+tmp[2747]*kernel[4]+tmp[2748]*kernel[5]+tmp[2846]*kernel[6]+tmp[2847]*kernel[7]+tmp[2848]*kernel[8];
				ans[2748]<=tmp[2647]*kernel[0]+tmp[2648]*kernel[1]+tmp[2649]*kernel[2]+tmp[2747]*kernel[3]+tmp[2748]*kernel[4]+tmp[2749]*kernel[5]+tmp[2847]*kernel[6]+tmp[2848]*kernel[7]+tmp[2849]*kernel[8];
				ans[2749]<=tmp[2648]*kernel[0]+tmp[2649]*kernel[1]+tmp[2650]*kernel[2]+tmp[2748]*kernel[3]+tmp[2749]*kernel[4]+tmp[2750]*kernel[5]+tmp[2848]*kernel[6]+tmp[2849]*kernel[7]+tmp[2850]*kernel[8];
				ans[2750]<=tmp[2649]*kernel[0]+tmp[2650]*kernel[1]+tmp[2651]*kernel[2]+tmp[2749]*kernel[3]+tmp[2750]*kernel[4]+tmp[2751]*kernel[5]+tmp[2849]*kernel[6]+tmp[2850]*kernel[7]+tmp[2851]*kernel[8];
				ans[2751]<=tmp[2650]*kernel[0]+tmp[2651]*kernel[1]+tmp[2652]*kernel[2]+tmp[2750]*kernel[3]+tmp[2751]*kernel[4]+tmp[2752]*kernel[5]+tmp[2850]*kernel[6]+tmp[2851]*kernel[7]+tmp[2852]*kernel[8];
				ans[2752]<=tmp[2651]*kernel[0]+tmp[2652]*kernel[1]+tmp[2653]*kernel[2]+tmp[2751]*kernel[3]+tmp[2752]*kernel[4]+tmp[2753]*kernel[5]+tmp[2851]*kernel[6]+tmp[2852]*kernel[7]+tmp[2853]*kernel[8];
				ans[2753]<=tmp[2652]*kernel[0]+tmp[2653]*kernel[1]+tmp[2654]*kernel[2]+tmp[2752]*kernel[3]+tmp[2753]*kernel[4]+tmp[2754]*kernel[5]+tmp[2852]*kernel[6]+tmp[2853]*kernel[7]+tmp[2854]*kernel[8];
				ans[2754]<=tmp[2653]*kernel[0]+tmp[2654]*kernel[1]+tmp[2655]*kernel[2]+tmp[2753]*kernel[3]+tmp[2754]*kernel[4]+tmp[2755]*kernel[5]+tmp[2853]*kernel[6]+tmp[2854]*kernel[7]+tmp[2855]*kernel[8];
				ans[2755]<=tmp[2654]*kernel[0]+tmp[2655]*kernel[1]+tmp[2656]*kernel[2]+tmp[2754]*kernel[3]+tmp[2755]*kernel[4]+tmp[2756]*kernel[5]+tmp[2854]*kernel[6]+tmp[2855]*kernel[7]+tmp[2856]*kernel[8];
				ans[2756]<=tmp[2655]*kernel[0]+tmp[2656]*kernel[1]+tmp[2657]*kernel[2]+tmp[2755]*kernel[3]+tmp[2756]*kernel[4]+tmp[2757]*kernel[5]+tmp[2855]*kernel[6]+tmp[2856]*kernel[7]+tmp[2857]*kernel[8];
				ans[2757]<=tmp[2656]*kernel[0]+tmp[2657]*kernel[1]+tmp[2658]*kernel[2]+tmp[2756]*kernel[3]+tmp[2757]*kernel[4]+tmp[2758]*kernel[5]+tmp[2856]*kernel[6]+tmp[2857]*kernel[7]+tmp[2858]*kernel[8];
				ans[2758]<=tmp[2657]*kernel[0]+tmp[2658]*kernel[1]+tmp[2659]*kernel[2]+tmp[2757]*kernel[3]+tmp[2758]*kernel[4]+tmp[2759]*kernel[5]+tmp[2857]*kernel[6]+tmp[2858]*kernel[7]+tmp[2859]*kernel[8];
				ans[2759]<=tmp[2658]*kernel[0]+tmp[2659]*kernel[1]+tmp[2660]*kernel[2]+tmp[2758]*kernel[3]+tmp[2759]*kernel[4]+tmp[2760]*kernel[5]+tmp[2858]*kernel[6]+tmp[2859]*kernel[7]+tmp[2860]*kernel[8];
				ans[2760]<=tmp[2659]*kernel[0]+tmp[2660]*kernel[1]+tmp[2661]*kernel[2]+tmp[2759]*kernel[3]+tmp[2760]*kernel[4]+tmp[2761]*kernel[5]+tmp[2859]*kernel[6]+tmp[2860]*kernel[7]+tmp[2861]*kernel[8];
				ans[2761]<=tmp[2660]*kernel[0]+tmp[2661]*kernel[1]+tmp[2662]*kernel[2]+tmp[2760]*kernel[3]+tmp[2761]*kernel[4]+tmp[2762]*kernel[5]+tmp[2860]*kernel[6]+tmp[2861]*kernel[7]+tmp[2862]*kernel[8];
				ans[2762]<=tmp[2661]*kernel[0]+tmp[2662]*kernel[1]+tmp[2663]*kernel[2]+tmp[2761]*kernel[3]+tmp[2762]*kernel[4]+tmp[2763]*kernel[5]+tmp[2861]*kernel[6]+tmp[2862]*kernel[7]+tmp[2863]*kernel[8];
				ans[2763]<=tmp[2662]*kernel[0]+tmp[2663]*kernel[1]+tmp[2664]*kernel[2]+tmp[2762]*kernel[3]+tmp[2763]*kernel[4]+tmp[2764]*kernel[5]+tmp[2862]*kernel[6]+tmp[2863]*kernel[7]+tmp[2864]*kernel[8];
				ans[2764]<=tmp[2663]*kernel[0]+tmp[2664]*kernel[1]+tmp[2665]*kernel[2]+tmp[2763]*kernel[3]+tmp[2764]*kernel[4]+tmp[2765]*kernel[5]+tmp[2863]*kernel[6]+tmp[2864]*kernel[7]+tmp[2865]*kernel[8];
				ans[2765]<=tmp[2664]*kernel[0]+tmp[2665]*kernel[1]+tmp[2666]*kernel[2]+tmp[2764]*kernel[3]+tmp[2765]*kernel[4]+tmp[2766]*kernel[5]+tmp[2864]*kernel[6]+tmp[2865]*kernel[7]+tmp[2866]*kernel[8];
				ans[2766]<=tmp[2665]*kernel[0]+tmp[2666]*kernel[1]+tmp[2667]*kernel[2]+tmp[2765]*kernel[3]+tmp[2766]*kernel[4]+tmp[2767]*kernel[5]+tmp[2865]*kernel[6]+tmp[2866]*kernel[7]+tmp[2867]*kernel[8];
				ans[2767]<=tmp[2666]*kernel[0]+tmp[2667]*kernel[1]+tmp[2668]*kernel[2]+tmp[2766]*kernel[3]+tmp[2767]*kernel[4]+tmp[2768]*kernel[5]+tmp[2866]*kernel[6]+tmp[2867]*kernel[7]+tmp[2868]*kernel[8];
				ans[2768]<=tmp[2667]*kernel[0]+tmp[2668]*kernel[1]+tmp[2669]*kernel[2]+tmp[2767]*kernel[3]+tmp[2768]*kernel[4]+tmp[2769]*kernel[5]+tmp[2867]*kernel[6]+tmp[2868]*kernel[7]+tmp[2869]*kernel[8];
				ans[2769]<=tmp[2668]*kernel[0]+tmp[2669]*kernel[1]+tmp[2670]*kernel[2]+tmp[2768]*kernel[3]+tmp[2769]*kernel[4]+tmp[2770]*kernel[5]+tmp[2868]*kernel[6]+tmp[2869]*kernel[7]+tmp[2870]*kernel[8];
				ans[2770]<=tmp[2669]*kernel[0]+tmp[2670]*kernel[1]+tmp[2671]*kernel[2]+tmp[2769]*kernel[3]+tmp[2770]*kernel[4]+tmp[2771]*kernel[5]+tmp[2869]*kernel[6]+tmp[2870]*kernel[7]+tmp[2871]*kernel[8];
				ans[2771]<=tmp[2670]*kernel[0]+tmp[2671]*kernel[1]+tmp[2672]*kernel[2]+tmp[2770]*kernel[3]+tmp[2771]*kernel[4]+tmp[2772]*kernel[5]+tmp[2870]*kernel[6]+tmp[2871]*kernel[7]+tmp[2872]*kernel[8];
				ans[2772]<=tmp[2671]*kernel[0]+tmp[2672]*kernel[1]+tmp[2673]*kernel[2]+tmp[2771]*kernel[3]+tmp[2772]*kernel[4]+tmp[2773]*kernel[5]+tmp[2871]*kernel[6]+tmp[2872]*kernel[7]+tmp[2873]*kernel[8];
				ans[2773]<=tmp[2672]*kernel[0]+tmp[2673]*kernel[1]+tmp[2674]*kernel[2]+tmp[2772]*kernel[3]+tmp[2773]*kernel[4]+tmp[2774]*kernel[5]+tmp[2872]*kernel[6]+tmp[2873]*kernel[7]+tmp[2874]*kernel[8];
				ans[2774]<=tmp[2673]*kernel[0]+tmp[2674]*kernel[1]+tmp[2675]*kernel[2]+tmp[2773]*kernel[3]+tmp[2774]*kernel[4]+tmp[2775]*kernel[5]+tmp[2873]*kernel[6]+tmp[2874]*kernel[7]+tmp[2875]*kernel[8];
				ans[2775]<=tmp[2674]*kernel[0]+tmp[2675]*kernel[1]+tmp[2676]*kernel[2]+tmp[2774]*kernel[3]+tmp[2775]*kernel[4]+tmp[2776]*kernel[5]+tmp[2874]*kernel[6]+tmp[2875]*kernel[7]+tmp[2876]*kernel[8];
				ans[2776]<=tmp[2675]*kernel[0]+tmp[2676]*kernel[1]+tmp[2677]*kernel[2]+tmp[2775]*kernel[3]+tmp[2776]*kernel[4]+tmp[2777]*kernel[5]+tmp[2875]*kernel[6]+tmp[2876]*kernel[7]+tmp[2877]*kernel[8];
				ans[2777]<=tmp[2676]*kernel[0]+tmp[2677]*kernel[1]+tmp[2678]*kernel[2]+tmp[2776]*kernel[3]+tmp[2777]*kernel[4]+tmp[2778]*kernel[5]+tmp[2876]*kernel[6]+tmp[2877]*kernel[7]+tmp[2878]*kernel[8];
				ans[2778]<=tmp[2677]*kernel[0]+tmp[2678]*kernel[1]+tmp[2679]*kernel[2]+tmp[2777]*kernel[3]+tmp[2778]*kernel[4]+tmp[2779]*kernel[5]+tmp[2877]*kernel[6]+tmp[2878]*kernel[7]+tmp[2879]*kernel[8];
				ans[2779]<=tmp[2678]*kernel[0]+tmp[2679]*kernel[1]+tmp[2680]*kernel[2]+tmp[2778]*kernel[3]+tmp[2779]*kernel[4]+tmp[2780]*kernel[5]+tmp[2878]*kernel[6]+tmp[2879]*kernel[7]+tmp[2880]*kernel[8];
				ans[2780]<=tmp[2679]*kernel[0]+tmp[2680]*kernel[1]+tmp[2681]*kernel[2]+tmp[2779]*kernel[3]+tmp[2780]*kernel[4]+tmp[2781]*kernel[5]+tmp[2879]*kernel[6]+tmp[2880]*kernel[7]+tmp[2881]*kernel[8];
				ans[2781]<=tmp[2680]*kernel[0]+tmp[2681]*kernel[1]+tmp[2682]*kernel[2]+tmp[2780]*kernel[3]+tmp[2781]*kernel[4]+tmp[2782]*kernel[5]+tmp[2880]*kernel[6]+tmp[2881]*kernel[7]+tmp[2882]*kernel[8];
				ans[2782]<=tmp[2681]*kernel[0]+tmp[2682]*kernel[1]+tmp[2683]*kernel[2]+tmp[2781]*kernel[3]+tmp[2782]*kernel[4]+tmp[2783]*kernel[5]+tmp[2881]*kernel[6]+tmp[2882]*kernel[7]+tmp[2883]*kernel[8];
				ans[2783]<=tmp[2682]*kernel[0]+tmp[2683]*kernel[1]+tmp[2684]*kernel[2]+tmp[2782]*kernel[3]+tmp[2783]*kernel[4]+tmp[2784]*kernel[5]+tmp[2882]*kernel[6]+tmp[2883]*kernel[7]+tmp[2884]*kernel[8];
				ans[2784]<=tmp[2683]*kernel[0]+tmp[2684]*kernel[1]+tmp[2685]*kernel[2]+tmp[2783]*kernel[3]+tmp[2784]*kernel[4]+tmp[2785]*kernel[5]+tmp[2883]*kernel[6]+tmp[2884]*kernel[7]+tmp[2885]*kernel[8];
				ans[2785]<=tmp[2684]*kernel[0]+tmp[2685]*kernel[1]+tmp[2686]*kernel[2]+tmp[2784]*kernel[3]+tmp[2785]*kernel[4]+tmp[2786]*kernel[5]+tmp[2884]*kernel[6]+tmp[2885]*kernel[7]+tmp[2886]*kernel[8];
				ans[2786]<=tmp[2685]*kernel[0]+tmp[2686]*kernel[1]+tmp[2687]*kernel[2]+tmp[2785]*kernel[3]+tmp[2786]*kernel[4]+tmp[2787]*kernel[5]+tmp[2885]*kernel[6]+tmp[2886]*kernel[7]+tmp[2887]*kernel[8];
				ans[2787]<=tmp[2686]*kernel[0]+tmp[2687]*kernel[1]+tmp[2688]*kernel[2]+tmp[2786]*kernel[3]+tmp[2787]*kernel[4]+tmp[2788]*kernel[5]+tmp[2886]*kernel[6]+tmp[2887]*kernel[7]+tmp[2888]*kernel[8];
				ans[2788]<=tmp[2687]*kernel[0]+tmp[2688]*kernel[1]+tmp[2689]*kernel[2]+tmp[2787]*kernel[3]+tmp[2788]*kernel[4]+tmp[2789]*kernel[5]+tmp[2887]*kernel[6]+tmp[2888]*kernel[7]+tmp[2889]*kernel[8];
				ans[2789]<=tmp[2688]*kernel[0]+tmp[2689]*kernel[1]+tmp[2690]*kernel[2]+tmp[2788]*kernel[3]+tmp[2789]*kernel[4]+tmp[2790]*kernel[5]+tmp[2888]*kernel[6]+tmp[2889]*kernel[7]+tmp[2890]*kernel[8];
				ans[2790]<=tmp[2689]*kernel[0]+tmp[2690]*kernel[1]+tmp[2691]*kernel[2]+tmp[2789]*kernel[3]+tmp[2790]*kernel[4]+tmp[2791]*kernel[5]+tmp[2889]*kernel[6]+tmp[2890]*kernel[7]+tmp[2891]*kernel[8];
				ans[2791]<=tmp[2690]*kernel[0]+tmp[2691]*kernel[1]+tmp[2692]*kernel[2]+tmp[2790]*kernel[3]+tmp[2791]*kernel[4]+tmp[2792]*kernel[5]+tmp[2890]*kernel[6]+tmp[2891]*kernel[7]+tmp[2892]*kernel[8];
				ans[2792]<=tmp[2691]*kernel[0]+tmp[2692]*kernel[1]+tmp[2693]*kernel[2]+tmp[2791]*kernel[3]+tmp[2792]*kernel[4]+tmp[2793]*kernel[5]+tmp[2891]*kernel[6]+tmp[2892]*kernel[7]+tmp[2893]*kernel[8];
				ans[2793]<=tmp[2692]*kernel[0]+tmp[2693]*kernel[1]+tmp[2694]*kernel[2]+tmp[2792]*kernel[3]+tmp[2793]*kernel[4]+tmp[2794]*kernel[5]+tmp[2892]*kernel[6]+tmp[2893]*kernel[7]+tmp[2894]*kernel[8];
				ans[2794]<=tmp[2693]*kernel[0]+tmp[2694]*kernel[1]+tmp[2695]*kernel[2]+tmp[2793]*kernel[3]+tmp[2794]*kernel[4]+tmp[2795]*kernel[5]+tmp[2893]*kernel[6]+tmp[2894]*kernel[7]+tmp[2895]*kernel[8];
				ans[2795]<=tmp[2694]*kernel[0]+tmp[2695]*kernel[1]+tmp[2696]*kernel[2]+tmp[2794]*kernel[3]+tmp[2795]*kernel[4]+tmp[2796]*kernel[5]+tmp[2894]*kernel[6]+tmp[2895]*kernel[7]+tmp[2896]*kernel[8];
				ans[2796]<=tmp[2695]*kernel[0]+tmp[2696]*kernel[1]+tmp[2697]*kernel[2]+tmp[2795]*kernel[3]+tmp[2796]*kernel[4]+tmp[2797]*kernel[5]+tmp[2895]*kernel[6]+tmp[2896]*kernel[7]+tmp[2897]*kernel[8];
				ans[2797]<=tmp[2696]*kernel[0]+tmp[2697]*kernel[1]+tmp[2698]*kernel[2]+tmp[2796]*kernel[3]+tmp[2797]*kernel[4]+tmp[2798]*kernel[5]+tmp[2896]*kernel[6]+tmp[2897]*kernel[7]+tmp[2898]*kernel[8];
				ans[2798]<=tmp[2697]*kernel[0]+tmp[2698]*kernel[1]+tmp[2699]*kernel[2]+tmp[2797]*kernel[3]+tmp[2798]*kernel[4]+tmp[2799]*kernel[5]+tmp[2897]*kernel[6]+tmp[2898]*kernel[7]+tmp[2899]*kernel[8];
				ans[2799]<=tmp[2698]*kernel[0]+tmp[2699]*kernel[1]+tmp[2798]*kernel[3]+tmp[2799]*kernel[4]+tmp[2898]*kernel[6]+tmp[2899]*kernel[7];
				ans[2800]<=tmp[2700]*kernel[1]+tmp[2701]*kernel[2]+tmp[2800]*kernel[4]+tmp[2801]*kernel[5]+tmp[2900]*kernel[7]+tmp[2901]*kernel[8];
				ans[2801]<=tmp[2700]*kernel[0]+tmp[2701]*kernel[1]+tmp[2702]*kernel[2]+tmp[2800]*kernel[3]+tmp[2801]*kernel[4]+tmp[2802]*kernel[5]+tmp[2900]*kernel[6]+tmp[2901]*kernel[7]+tmp[2902]*kernel[8];
				ans[2802]<=tmp[2701]*kernel[0]+tmp[2702]*kernel[1]+tmp[2703]*kernel[2]+tmp[2801]*kernel[3]+tmp[2802]*kernel[4]+tmp[2803]*kernel[5]+tmp[2901]*kernel[6]+tmp[2902]*kernel[7]+tmp[2903]*kernel[8];
				ans[2803]<=tmp[2702]*kernel[0]+tmp[2703]*kernel[1]+tmp[2704]*kernel[2]+tmp[2802]*kernel[3]+tmp[2803]*kernel[4]+tmp[2804]*kernel[5]+tmp[2902]*kernel[6]+tmp[2903]*kernel[7]+tmp[2904]*kernel[8];
				ans[2804]<=tmp[2703]*kernel[0]+tmp[2704]*kernel[1]+tmp[2705]*kernel[2]+tmp[2803]*kernel[3]+tmp[2804]*kernel[4]+tmp[2805]*kernel[5]+tmp[2903]*kernel[6]+tmp[2904]*kernel[7]+tmp[2905]*kernel[8];
				ans[2805]<=tmp[2704]*kernel[0]+tmp[2705]*kernel[1]+tmp[2706]*kernel[2]+tmp[2804]*kernel[3]+tmp[2805]*kernel[4]+tmp[2806]*kernel[5]+tmp[2904]*kernel[6]+tmp[2905]*kernel[7]+tmp[2906]*kernel[8];
				ans[2806]<=tmp[2705]*kernel[0]+tmp[2706]*kernel[1]+tmp[2707]*kernel[2]+tmp[2805]*kernel[3]+tmp[2806]*kernel[4]+tmp[2807]*kernel[5]+tmp[2905]*kernel[6]+tmp[2906]*kernel[7]+tmp[2907]*kernel[8];
				ans[2807]<=tmp[2706]*kernel[0]+tmp[2707]*kernel[1]+tmp[2708]*kernel[2]+tmp[2806]*kernel[3]+tmp[2807]*kernel[4]+tmp[2808]*kernel[5]+tmp[2906]*kernel[6]+tmp[2907]*kernel[7]+tmp[2908]*kernel[8];
				ans[2808]<=tmp[2707]*kernel[0]+tmp[2708]*kernel[1]+tmp[2709]*kernel[2]+tmp[2807]*kernel[3]+tmp[2808]*kernel[4]+tmp[2809]*kernel[5]+tmp[2907]*kernel[6]+tmp[2908]*kernel[7]+tmp[2909]*kernel[8];
				ans[2809]<=tmp[2708]*kernel[0]+tmp[2709]*kernel[1]+tmp[2710]*kernel[2]+tmp[2808]*kernel[3]+tmp[2809]*kernel[4]+tmp[2810]*kernel[5]+tmp[2908]*kernel[6]+tmp[2909]*kernel[7]+tmp[2910]*kernel[8];
				ans[2810]<=tmp[2709]*kernel[0]+tmp[2710]*kernel[1]+tmp[2711]*kernel[2]+tmp[2809]*kernel[3]+tmp[2810]*kernel[4]+tmp[2811]*kernel[5]+tmp[2909]*kernel[6]+tmp[2910]*kernel[7]+tmp[2911]*kernel[8];
				ans[2811]<=tmp[2710]*kernel[0]+tmp[2711]*kernel[1]+tmp[2712]*kernel[2]+tmp[2810]*kernel[3]+tmp[2811]*kernel[4]+tmp[2812]*kernel[5]+tmp[2910]*kernel[6]+tmp[2911]*kernel[7]+tmp[2912]*kernel[8];
				ans[2812]<=tmp[2711]*kernel[0]+tmp[2712]*kernel[1]+tmp[2713]*kernel[2]+tmp[2811]*kernel[3]+tmp[2812]*kernel[4]+tmp[2813]*kernel[5]+tmp[2911]*kernel[6]+tmp[2912]*kernel[7]+tmp[2913]*kernel[8];
				ans[2813]<=tmp[2712]*kernel[0]+tmp[2713]*kernel[1]+tmp[2714]*kernel[2]+tmp[2812]*kernel[3]+tmp[2813]*kernel[4]+tmp[2814]*kernel[5]+tmp[2912]*kernel[6]+tmp[2913]*kernel[7]+tmp[2914]*kernel[8];
				ans[2814]<=tmp[2713]*kernel[0]+tmp[2714]*kernel[1]+tmp[2715]*kernel[2]+tmp[2813]*kernel[3]+tmp[2814]*kernel[4]+tmp[2815]*kernel[5]+tmp[2913]*kernel[6]+tmp[2914]*kernel[7]+tmp[2915]*kernel[8];
				ans[2815]<=tmp[2714]*kernel[0]+tmp[2715]*kernel[1]+tmp[2716]*kernel[2]+tmp[2814]*kernel[3]+tmp[2815]*kernel[4]+tmp[2816]*kernel[5]+tmp[2914]*kernel[6]+tmp[2915]*kernel[7]+tmp[2916]*kernel[8];
				ans[2816]<=tmp[2715]*kernel[0]+tmp[2716]*kernel[1]+tmp[2717]*kernel[2]+tmp[2815]*kernel[3]+tmp[2816]*kernel[4]+tmp[2817]*kernel[5]+tmp[2915]*kernel[6]+tmp[2916]*kernel[7]+tmp[2917]*kernel[8];
				ans[2817]<=tmp[2716]*kernel[0]+tmp[2717]*kernel[1]+tmp[2718]*kernel[2]+tmp[2816]*kernel[3]+tmp[2817]*kernel[4]+tmp[2818]*kernel[5]+tmp[2916]*kernel[6]+tmp[2917]*kernel[7]+tmp[2918]*kernel[8];
				ans[2818]<=tmp[2717]*kernel[0]+tmp[2718]*kernel[1]+tmp[2719]*kernel[2]+tmp[2817]*kernel[3]+tmp[2818]*kernel[4]+tmp[2819]*kernel[5]+tmp[2917]*kernel[6]+tmp[2918]*kernel[7]+tmp[2919]*kernel[8];
				ans[2819]<=tmp[2718]*kernel[0]+tmp[2719]*kernel[1]+tmp[2720]*kernel[2]+tmp[2818]*kernel[3]+tmp[2819]*kernel[4]+tmp[2820]*kernel[5]+tmp[2918]*kernel[6]+tmp[2919]*kernel[7]+tmp[2920]*kernel[8];
				ans[2820]<=tmp[2719]*kernel[0]+tmp[2720]*kernel[1]+tmp[2721]*kernel[2]+tmp[2819]*kernel[3]+tmp[2820]*kernel[4]+tmp[2821]*kernel[5]+tmp[2919]*kernel[6]+tmp[2920]*kernel[7]+tmp[2921]*kernel[8];
				ans[2821]<=tmp[2720]*kernel[0]+tmp[2721]*kernel[1]+tmp[2722]*kernel[2]+tmp[2820]*kernel[3]+tmp[2821]*kernel[4]+tmp[2822]*kernel[5]+tmp[2920]*kernel[6]+tmp[2921]*kernel[7]+tmp[2922]*kernel[8];
				ans[2822]<=tmp[2721]*kernel[0]+tmp[2722]*kernel[1]+tmp[2723]*kernel[2]+tmp[2821]*kernel[3]+tmp[2822]*kernel[4]+tmp[2823]*kernel[5]+tmp[2921]*kernel[6]+tmp[2922]*kernel[7]+tmp[2923]*kernel[8];
				ans[2823]<=tmp[2722]*kernel[0]+tmp[2723]*kernel[1]+tmp[2724]*kernel[2]+tmp[2822]*kernel[3]+tmp[2823]*kernel[4]+tmp[2824]*kernel[5]+tmp[2922]*kernel[6]+tmp[2923]*kernel[7]+tmp[2924]*kernel[8];
				ans[2824]<=tmp[2723]*kernel[0]+tmp[2724]*kernel[1]+tmp[2725]*kernel[2]+tmp[2823]*kernel[3]+tmp[2824]*kernel[4]+tmp[2825]*kernel[5]+tmp[2923]*kernel[6]+tmp[2924]*kernel[7]+tmp[2925]*kernel[8];
				ans[2825]<=tmp[2724]*kernel[0]+tmp[2725]*kernel[1]+tmp[2726]*kernel[2]+tmp[2824]*kernel[3]+tmp[2825]*kernel[4]+tmp[2826]*kernel[5]+tmp[2924]*kernel[6]+tmp[2925]*kernel[7]+tmp[2926]*kernel[8];
				ans[2826]<=tmp[2725]*kernel[0]+tmp[2726]*kernel[1]+tmp[2727]*kernel[2]+tmp[2825]*kernel[3]+tmp[2826]*kernel[4]+tmp[2827]*kernel[5]+tmp[2925]*kernel[6]+tmp[2926]*kernel[7]+tmp[2927]*kernel[8];
				ans[2827]<=tmp[2726]*kernel[0]+tmp[2727]*kernel[1]+tmp[2728]*kernel[2]+tmp[2826]*kernel[3]+tmp[2827]*kernel[4]+tmp[2828]*kernel[5]+tmp[2926]*kernel[6]+tmp[2927]*kernel[7]+tmp[2928]*kernel[8];
				ans[2828]<=tmp[2727]*kernel[0]+tmp[2728]*kernel[1]+tmp[2729]*kernel[2]+tmp[2827]*kernel[3]+tmp[2828]*kernel[4]+tmp[2829]*kernel[5]+tmp[2927]*kernel[6]+tmp[2928]*kernel[7]+tmp[2929]*kernel[8];
				ans[2829]<=tmp[2728]*kernel[0]+tmp[2729]*kernel[1]+tmp[2730]*kernel[2]+tmp[2828]*kernel[3]+tmp[2829]*kernel[4]+tmp[2830]*kernel[5]+tmp[2928]*kernel[6]+tmp[2929]*kernel[7]+tmp[2930]*kernel[8];
				ans[2830]<=tmp[2729]*kernel[0]+tmp[2730]*kernel[1]+tmp[2731]*kernel[2]+tmp[2829]*kernel[3]+tmp[2830]*kernel[4]+tmp[2831]*kernel[5]+tmp[2929]*kernel[6]+tmp[2930]*kernel[7]+tmp[2931]*kernel[8];
				ans[2831]<=tmp[2730]*kernel[0]+tmp[2731]*kernel[1]+tmp[2732]*kernel[2]+tmp[2830]*kernel[3]+tmp[2831]*kernel[4]+tmp[2832]*kernel[5]+tmp[2930]*kernel[6]+tmp[2931]*kernel[7]+tmp[2932]*kernel[8];
				ans[2832]<=tmp[2731]*kernel[0]+tmp[2732]*kernel[1]+tmp[2733]*kernel[2]+tmp[2831]*kernel[3]+tmp[2832]*kernel[4]+tmp[2833]*kernel[5]+tmp[2931]*kernel[6]+tmp[2932]*kernel[7]+tmp[2933]*kernel[8];
				ans[2833]<=tmp[2732]*kernel[0]+tmp[2733]*kernel[1]+tmp[2734]*kernel[2]+tmp[2832]*kernel[3]+tmp[2833]*kernel[4]+tmp[2834]*kernel[5]+tmp[2932]*kernel[6]+tmp[2933]*kernel[7]+tmp[2934]*kernel[8];
				ans[2834]<=tmp[2733]*kernel[0]+tmp[2734]*kernel[1]+tmp[2735]*kernel[2]+tmp[2833]*kernel[3]+tmp[2834]*kernel[4]+tmp[2835]*kernel[5]+tmp[2933]*kernel[6]+tmp[2934]*kernel[7]+tmp[2935]*kernel[8];
				ans[2835]<=tmp[2734]*kernel[0]+tmp[2735]*kernel[1]+tmp[2736]*kernel[2]+tmp[2834]*kernel[3]+tmp[2835]*kernel[4]+tmp[2836]*kernel[5]+tmp[2934]*kernel[6]+tmp[2935]*kernel[7]+tmp[2936]*kernel[8];
				ans[2836]<=tmp[2735]*kernel[0]+tmp[2736]*kernel[1]+tmp[2737]*kernel[2]+tmp[2835]*kernel[3]+tmp[2836]*kernel[4]+tmp[2837]*kernel[5]+tmp[2935]*kernel[6]+tmp[2936]*kernel[7]+tmp[2937]*kernel[8];
				ans[2837]<=tmp[2736]*kernel[0]+tmp[2737]*kernel[1]+tmp[2738]*kernel[2]+tmp[2836]*kernel[3]+tmp[2837]*kernel[4]+tmp[2838]*kernel[5]+tmp[2936]*kernel[6]+tmp[2937]*kernel[7]+tmp[2938]*kernel[8];
				ans[2838]<=tmp[2737]*kernel[0]+tmp[2738]*kernel[1]+tmp[2739]*kernel[2]+tmp[2837]*kernel[3]+tmp[2838]*kernel[4]+tmp[2839]*kernel[5]+tmp[2937]*kernel[6]+tmp[2938]*kernel[7]+tmp[2939]*kernel[8];
				ans[2839]<=tmp[2738]*kernel[0]+tmp[2739]*kernel[1]+tmp[2740]*kernel[2]+tmp[2838]*kernel[3]+tmp[2839]*kernel[4]+tmp[2840]*kernel[5]+tmp[2938]*kernel[6]+tmp[2939]*kernel[7]+tmp[2940]*kernel[8];
				ans[2840]<=tmp[2739]*kernel[0]+tmp[2740]*kernel[1]+tmp[2741]*kernel[2]+tmp[2839]*kernel[3]+tmp[2840]*kernel[4]+tmp[2841]*kernel[5]+tmp[2939]*kernel[6]+tmp[2940]*kernel[7]+tmp[2941]*kernel[8];
				ans[2841]<=tmp[2740]*kernel[0]+tmp[2741]*kernel[1]+tmp[2742]*kernel[2]+tmp[2840]*kernel[3]+tmp[2841]*kernel[4]+tmp[2842]*kernel[5]+tmp[2940]*kernel[6]+tmp[2941]*kernel[7]+tmp[2942]*kernel[8];
				ans[2842]<=tmp[2741]*kernel[0]+tmp[2742]*kernel[1]+tmp[2743]*kernel[2]+tmp[2841]*kernel[3]+tmp[2842]*kernel[4]+tmp[2843]*kernel[5]+tmp[2941]*kernel[6]+tmp[2942]*kernel[7]+tmp[2943]*kernel[8];
				ans[2843]<=tmp[2742]*kernel[0]+tmp[2743]*kernel[1]+tmp[2744]*kernel[2]+tmp[2842]*kernel[3]+tmp[2843]*kernel[4]+tmp[2844]*kernel[5]+tmp[2942]*kernel[6]+tmp[2943]*kernel[7]+tmp[2944]*kernel[8];
				ans[2844]<=tmp[2743]*kernel[0]+tmp[2744]*kernel[1]+tmp[2745]*kernel[2]+tmp[2843]*kernel[3]+tmp[2844]*kernel[4]+tmp[2845]*kernel[5]+tmp[2943]*kernel[6]+tmp[2944]*kernel[7]+tmp[2945]*kernel[8];
				ans[2845]<=tmp[2744]*kernel[0]+tmp[2745]*kernel[1]+tmp[2746]*kernel[2]+tmp[2844]*kernel[3]+tmp[2845]*kernel[4]+tmp[2846]*kernel[5]+tmp[2944]*kernel[6]+tmp[2945]*kernel[7]+tmp[2946]*kernel[8];
				ans[2846]<=tmp[2745]*kernel[0]+tmp[2746]*kernel[1]+tmp[2747]*kernel[2]+tmp[2845]*kernel[3]+tmp[2846]*kernel[4]+tmp[2847]*kernel[5]+tmp[2945]*kernel[6]+tmp[2946]*kernel[7]+tmp[2947]*kernel[8];
				ans[2847]<=tmp[2746]*kernel[0]+tmp[2747]*kernel[1]+tmp[2748]*kernel[2]+tmp[2846]*kernel[3]+tmp[2847]*kernel[4]+tmp[2848]*kernel[5]+tmp[2946]*kernel[6]+tmp[2947]*kernel[7]+tmp[2948]*kernel[8];
				ans[2848]<=tmp[2747]*kernel[0]+tmp[2748]*kernel[1]+tmp[2749]*kernel[2]+tmp[2847]*kernel[3]+tmp[2848]*kernel[4]+tmp[2849]*kernel[5]+tmp[2947]*kernel[6]+tmp[2948]*kernel[7]+tmp[2949]*kernel[8];
				ans[2849]<=tmp[2748]*kernel[0]+tmp[2749]*kernel[1]+tmp[2750]*kernel[2]+tmp[2848]*kernel[3]+tmp[2849]*kernel[4]+tmp[2850]*kernel[5]+tmp[2948]*kernel[6]+tmp[2949]*kernel[7]+tmp[2950]*kernel[8];
				ans[2850]<=tmp[2749]*kernel[0]+tmp[2750]*kernel[1]+tmp[2751]*kernel[2]+tmp[2849]*kernel[3]+tmp[2850]*kernel[4]+tmp[2851]*kernel[5]+tmp[2949]*kernel[6]+tmp[2950]*kernel[7]+tmp[2951]*kernel[8];
				ans[2851]<=tmp[2750]*kernel[0]+tmp[2751]*kernel[1]+tmp[2752]*kernel[2]+tmp[2850]*kernel[3]+tmp[2851]*kernel[4]+tmp[2852]*kernel[5]+tmp[2950]*kernel[6]+tmp[2951]*kernel[7]+tmp[2952]*kernel[8];
				ans[2852]<=tmp[2751]*kernel[0]+tmp[2752]*kernel[1]+tmp[2753]*kernel[2]+tmp[2851]*kernel[3]+tmp[2852]*kernel[4]+tmp[2853]*kernel[5]+tmp[2951]*kernel[6]+tmp[2952]*kernel[7]+tmp[2953]*kernel[8];
				ans[2853]<=tmp[2752]*kernel[0]+tmp[2753]*kernel[1]+tmp[2754]*kernel[2]+tmp[2852]*kernel[3]+tmp[2853]*kernel[4]+tmp[2854]*kernel[5]+tmp[2952]*kernel[6]+tmp[2953]*kernel[7]+tmp[2954]*kernel[8];
				ans[2854]<=tmp[2753]*kernel[0]+tmp[2754]*kernel[1]+tmp[2755]*kernel[2]+tmp[2853]*kernel[3]+tmp[2854]*kernel[4]+tmp[2855]*kernel[5]+tmp[2953]*kernel[6]+tmp[2954]*kernel[7]+tmp[2955]*kernel[8];
				ans[2855]<=tmp[2754]*kernel[0]+tmp[2755]*kernel[1]+tmp[2756]*kernel[2]+tmp[2854]*kernel[3]+tmp[2855]*kernel[4]+tmp[2856]*kernel[5]+tmp[2954]*kernel[6]+tmp[2955]*kernel[7]+tmp[2956]*kernel[8];
				ans[2856]<=tmp[2755]*kernel[0]+tmp[2756]*kernel[1]+tmp[2757]*kernel[2]+tmp[2855]*kernel[3]+tmp[2856]*kernel[4]+tmp[2857]*kernel[5]+tmp[2955]*kernel[6]+tmp[2956]*kernel[7]+tmp[2957]*kernel[8];
				ans[2857]<=tmp[2756]*kernel[0]+tmp[2757]*kernel[1]+tmp[2758]*kernel[2]+tmp[2856]*kernel[3]+tmp[2857]*kernel[4]+tmp[2858]*kernel[5]+tmp[2956]*kernel[6]+tmp[2957]*kernel[7]+tmp[2958]*kernel[8];
				ans[2858]<=tmp[2757]*kernel[0]+tmp[2758]*kernel[1]+tmp[2759]*kernel[2]+tmp[2857]*kernel[3]+tmp[2858]*kernel[4]+tmp[2859]*kernel[5]+tmp[2957]*kernel[6]+tmp[2958]*kernel[7]+tmp[2959]*kernel[8];
				ans[2859]<=tmp[2758]*kernel[0]+tmp[2759]*kernel[1]+tmp[2760]*kernel[2]+tmp[2858]*kernel[3]+tmp[2859]*kernel[4]+tmp[2860]*kernel[5]+tmp[2958]*kernel[6]+tmp[2959]*kernel[7]+tmp[2960]*kernel[8];
				ans[2860]<=tmp[2759]*kernel[0]+tmp[2760]*kernel[1]+tmp[2761]*kernel[2]+tmp[2859]*kernel[3]+tmp[2860]*kernel[4]+tmp[2861]*kernel[5]+tmp[2959]*kernel[6]+tmp[2960]*kernel[7]+tmp[2961]*kernel[8];
				ans[2861]<=tmp[2760]*kernel[0]+tmp[2761]*kernel[1]+tmp[2762]*kernel[2]+tmp[2860]*kernel[3]+tmp[2861]*kernel[4]+tmp[2862]*kernel[5]+tmp[2960]*kernel[6]+tmp[2961]*kernel[7]+tmp[2962]*kernel[8];
				ans[2862]<=tmp[2761]*kernel[0]+tmp[2762]*kernel[1]+tmp[2763]*kernel[2]+tmp[2861]*kernel[3]+tmp[2862]*kernel[4]+tmp[2863]*kernel[5]+tmp[2961]*kernel[6]+tmp[2962]*kernel[7]+tmp[2963]*kernel[8];
				ans[2863]<=tmp[2762]*kernel[0]+tmp[2763]*kernel[1]+tmp[2764]*kernel[2]+tmp[2862]*kernel[3]+tmp[2863]*kernel[4]+tmp[2864]*kernel[5]+tmp[2962]*kernel[6]+tmp[2963]*kernel[7]+tmp[2964]*kernel[8];
				ans[2864]<=tmp[2763]*kernel[0]+tmp[2764]*kernel[1]+tmp[2765]*kernel[2]+tmp[2863]*kernel[3]+tmp[2864]*kernel[4]+tmp[2865]*kernel[5]+tmp[2963]*kernel[6]+tmp[2964]*kernel[7]+tmp[2965]*kernel[8];
				ans[2865]<=tmp[2764]*kernel[0]+tmp[2765]*kernel[1]+tmp[2766]*kernel[2]+tmp[2864]*kernel[3]+tmp[2865]*kernel[4]+tmp[2866]*kernel[5]+tmp[2964]*kernel[6]+tmp[2965]*kernel[7]+tmp[2966]*kernel[8];
				ans[2866]<=tmp[2765]*kernel[0]+tmp[2766]*kernel[1]+tmp[2767]*kernel[2]+tmp[2865]*kernel[3]+tmp[2866]*kernel[4]+tmp[2867]*kernel[5]+tmp[2965]*kernel[6]+tmp[2966]*kernel[7]+tmp[2967]*kernel[8];
				ans[2867]<=tmp[2766]*kernel[0]+tmp[2767]*kernel[1]+tmp[2768]*kernel[2]+tmp[2866]*kernel[3]+tmp[2867]*kernel[4]+tmp[2868]*kernel[5]+tmp[2966]*kernel[6]+tmp[2967]*kernel[7]+tmp[2968]*kernel[8];
				ans[2868]<=tmp[2767]*kernel[0]+tmp[2768]*kernel[1]+tmp[2769]*kernel[2]+tmp[2867]*kernel[3]+tmp[2868]*kernel[4]+tmp[2869]*kernel[5]+tmp[2967]*kernel[6]+tmp[2968]*kernel[7]+tmp[2969]*kernel[8];
				ans[2869]<=tmp[2768]*kernel[0]+tmp[2769]*kernel[1]+tmp[2770]*kernel[2]+tmp[2868]*kernel[3]+tmp[2869]*kernel[4]+tmp[2870]*kernel[5]+tmp[2968]*kernel[6]+tmp[2969]*kernel[7]+tmp[2970]*kernel[8];
				ans[2870]<=tmp[2769]*kernel[0]+tmp[2770]*kernel[1]+tmp[2771]*kernel[2]+tmp[2869]*kernel[3]+tmp[2870]*kernel[4]+tmp[2871]*kernel[5]+tmp[2969]*kernel[6]+tmp[2970]*kernel[7]+tmp[2971]*kernel[8];
				ans[2871]<=tmp[2770]*kernel[0]+tmp[2771]*kernel[1]+tmp[2772]*kernel[2]+tmp[2870]*kernel[3]+tmp[2871]*kernel[4]+tmp[2872]*kernel[5]+tmp[2970]*kernel[6]+tmp[2971]*kernel[7]+tmp[2972]*kernel[8];
				ans[2872]<=tmp[2771]*kernel[0]+tmp[2772]*kernel[1]+tmp[2773]*kernel[2]+tmp[2871]*kernel[3]+tmp[2872]*kernel[4]+tmp[2873]*kernel[5]+tmp[2971]*kernel[6]+tmp[2972]*kernel[7]+tmp[2973]*kernel[8];
				ans[2873]<=tmp[2772]*kernel[0]+tmp[2773]*kernel[1]+tmp[2774]*kernel[2]+tmp[2872]*kernel[3]+tmp[2873]*kernel[4]+tmp[2874]*kernel[5]+tmp[2972]*kernel[6]+tmp[2973]*kernel[7]+tmp[2974]*kernel[8];
				ans[2874]<=tmp[2773]*kernel[0]+tmp[2774]*kernel[1]+tmp[2775]*kernel[2]+tmp[2873]*kernel[3]+tmp[2874]*kernel[4]+tmp[2875]*kernel[5]+tmp[2973]*kernel[6]+tmp[2974]*kernel[7]+tmp[2975]*kernel[8];
				ans[2875]<=tmp[2774]*kernel[0]+tmp[2775]*kernel[1]+tmp[2776]*kernel[2]+tmp[2874]*kernel[3]+tmp[2875]*kernel[4]+tmp[2876]*kernel[5]+tmp[2974]*kernel[6]+tmp[2975]*kernel[7]+tmp[2976]*kernel[8];
				ans[2876]<=tmp[2775]*kernel[0]+tmp[2776]*kernel[1]+tmp[2777]*kernel[2]+tmp[2875]*kernel[3]+tmp[2876]*kernel[4]+tmp[2877]*kernel[5]+tmp[2975]*kernel[6]+tmp[2976]*kernel[7]+tmp[2977]*kernel[8];
				ans[2877]<=tmp[2776]*kernel[0]+tmp[2777]*kernel[1]+tmp[2778]*kernel[2]+tmp[2876]*kernel[3]+tmp[2877]*kernel[4]+tmp[2878]*kernel[5]+tmp[2976]*kernel[6]+tmp[2977]*kernel[7]+tmp[2978]*kernel[8];
				ans[2878]<=tmp[2777]*kernel[0]+tmp[2778]*kernel[1]+tmp[2779]*kernel[2]+tmp[2877]*kernel[3]+tmp[2878]*kernel[4]+tmp[2879]*kernel[5]+tmp[2977]*kernel[6]+tmp[2978]*kernel[7]+tmp[2979]*kernel[8];
				ans[2879]<=tmp[2778]*kernel[0]+tmp[2779]*kernel[1]+tmp[2780]*kernel[2]+tmp[2878]*kernel[3]+tmp[2879]*kernel[4]+tmp[2880]*kernel[5]+tmp[2978]*kernel[6]+tmp[2979]*kernel[7]+tmp[2980]*kernel[8];
				ans[2880]<=tmp[2779]*kernel[0]+tmp[2780]*kernel[1]+tmp[2781]*kernel[2]+tmp[2879]*kernel[3]+tmp[2880]*kernel[4]+tmp[2881]*kernel[5]+tmp[2979]*kernel[6]+tmp[2980]*kernel[7]+tmp[2981]*kernel[8];
				ans[2881]<=tmp[2780]*kernel[0]+tmp[2781]*kernel[1]+tmp[2782]*kernel[2]+tmp[2880]*kernel[3]+tmp[2881]*kernel[4]+tmp[2882]*kernel[5]+tmp[2980]*kernel[6]+tmp[2981]*kernel[7]+tmp[2982]*kernel[8];
				ans[2882]<=tmp[2781]*kernel[0]+tmp[2782]*kernel[1]+tmp[2783]*kernel[2]+tmp[2881]*kernel[3]+tmp[2882]*kernel[4]+tmp[2883]*kernel[5]+tmp[2981]*kernel[6]+tmp[2982]*kernel[7]+tmp[2983]*kernel[8];
				ans[2883]<=tmp[2782]*kernel[0]+tmp[2783]*kernel[1]+tmp[2784]*kernel[2]+tmp[2882]*kernel[3]+tmp[2883]*kernel[4]+tmp[2884]*kernel[5]+tmp[2982]*kernel[6]+tmp[2983]*kernel[7]+tmp[2984]*kernel[8];
				ans[2884]<=tmp[2783]*kernel[0]+tmp[2784]*kernel[1]+tmp[2785]*kernel[2]+tmp[2883]*kernel[3]+tmp[2884]*kernel[4]+tmp[2885]*kernel[5]+tmp[2983]*kernel[6]+tmp[2984]*kernel[7]+tmp[2985]*kernel[8];
				ans[2885]<=tmp[2784]*kernel[0]+tmp[2785]*kernel[1]+tmp[2786]*kernel[2]+tmp[2884]*kernel[3]+tmp[2885]*kernel[4]+tmp[2886]*kernel[5]+tmp[2984]*kernel[6]+tmp[2985]*kernel[7]+tmp[2986]*kernel[8];
				ans[2886]<=tmp[2785]*kernel[0]+tmp[2786]*kernel[1]+tmp[2787]*kernel[2]+tmp[2885]*kernel[3]+tmp[2886]*kernel[4]+tmp[2887]*kernel[5]+tmp[2985]*kernel[6]+tmp[2986]*kernel[7]+tmp[2987]*kernel[8];
				ans[2887]<=tmp[2786]*kernel[0]+tmp[2787]*kernel[1]+tmp[2788]*kernel[2]+tmp[2886]*kernel[3]+tmp[2887]*kernel[4]+tmp[2888]*kernel[5]+tmp[2986]*kernel[6]+tmp[2987]*kernel[7]+tmp[2988]*kernel[8];
				ans[2888]<=tmp[2787]*kernel[0]+tmp[2788]*kernel[1]+tmp[2789]*kernel[2]+tmp[2887]*kernel[3]+tmp[2888]*kernel[4]+tmp[2889]*kernel[5]+tmp[2987]*kernel[6]+tmp[2988]*kernel[7]+tmp[2989]*kernel[8];
				ans[2889]<=tmp[2788]*kernel[0]+tmp[2789]*kernel[1]+tmp[2790]*kernel[2]+tmp[2888]*kernel[3]+tmp[2889]*kernel[4]+tmp[2890]*kernel[5]+tmp[2988]*kernel[6]+tmp[2989]*kernel[7]+tmp[2990]*kernel[8];
				ans[2890]<=tmp[2789]*kernel[0]+tmp[2790]*kernel[1]+tmp[2791]*kernel[2]+tmp[2889]*kernel[3]+tmp[2890]*kernel[4]+tmp[2891]*kernel[5]+tmp[2989]*kernel[6]+tmp[2990]*kernel[7]+tmp[2991]*kernel[8];
				ans[2891]<=tmp[2790]*kernel[0]+tmp[2791]*kernel[1]+tmp[2792]*kernel[2]+tmp[2890]*kernel[3]+tmp[2891]*kernel[4]+tmp[2892]*kernel[5]+tmp[2990]*kernel[6]+tmp[2991]*kernel[7]+tmp[2992]*kernel[8];
				ans[2892]<=tmp[2791]*kernel[0]+tmp[2792]*kernel[1]+tmp[2793]*kernel[2]+tmp[2891]*kernel[3]+tmp[2892]*kernel[4]+tmp[2893]*kernel[5]+tmp[2991]*kernel[6]+tmp[2992]*kernel[7]+tmp[2993]*kernel[8];
				ans[2893]<=tmp[2792]*kernel[0]+tmp[2793]*kernel[1]+tmp[2794]*kernel[2]+tmp[2892]*kernel[3]+tmp[2893]*kernel[4]+tmp[2894]*kernel[5]+tmp[2992]*kernel[6]+tmp[2993]*kernel[7]+tmp[2994]*kernel[8];
				ans[2894]<=tmp[2793]*kernel[0]+tmp[2794]*kernel[1]+tmp[2795]*kernel[2]+tmp[2893]*kernel[3]+tmp[2894]*kernel[4]+tmp[2895]*kernel[5]+tmp[2993]*kernel[6]+tmp[2994]*kernel[7]+tmp[2995]*kernel[8];
				ans[2895]<=tmp[2794]*kernel[0]+tmp[2795]*kernel[1]+tmp[2796]*kernel[2]+tmp[2894]*kernel[3]+tmp[2895]*kernel[4]+tmp[2896]*kernel[5]+tmp[2994]*kernel[6]+tmp[2995]*kernel[7]+tmp[2996]*kernel[8];
				ans[2896]<=tmp[2795]*kernel[0]+tmp[2796]*kernel[1]+tmp[2797]*kernel[2]+tmp[2895]*kernel[3]+tmp[2896]*kernel[4]+tmp[2897]*kernel[5]+tmp[2995]*kernel[6]+tmp[2996]*kernel[7]+tmp[2997]*kernel[8];
				ans[2897]<=tmp[2796]*kernel[0]+tmp[2797]*kernel[1]+tmp[2798]*kernel[2]+tmp[2896]*kernel[3]+tmp[2897]*kernel[4]+tmp[2898]*kernel[5]+tmp[2996]*kernel[6]+tmp[2997]*kernel[7]+tmp[2998]*kernel[8];
				ans[2898]<=tmp[2797]*kernel[0]+tmp[2798]*kernel[1]+tmp[2799]*kernel[2]+tmp[2897]*kernel[3]+tmp[2898]*kernel[4]+tmp[2899]*kernel[5]+tmp[2997]*kernel[6]+tmp[2998]*kernel[7]+tmp[2999]*kernel[8];
				ans[2899]<=tmp[2798]*kernel[0]+tmp[2799]*kernel[1]+tmp[2898]*kernel[3]+tmp[2899]*kernel[4]+tmp[2998]*kernel[6]+tmp[2999]*kernel[7];
				ans[2900]<=tmp[2800]*kernel[1]+tmp[2801]*kernel[2]+tmp[2900]*kernel[4]+tmp[2901]*kernel[5]+tmp[3000]*kernel[7]+tmp[3001]*kernel[8];
				ans[2901]<=tmp[2800]*kernel[0]+tmp[2801]*kernel[1]+tmp[2802]*kernel[2]+tmp[2900]*kernel[3]+tmp[2901]*kernel[4]+tmp[2902]*kernel[5]+tmp[3000]*kernel[6]+tmp[3001]*kernel[7]+tmp[3002]*kernel[8];
				ans[2902]<=tmp[2801]*kernel[0]+tmp[2802]*kernel[1]+tmp[2803]*kernel[2]+tmp[2901]*kernel[3]+tmp[2902]*kernel[4]+tmp[2903]*kernel[5]+tmp[3001]*kernel[6]+tmp[3002]*kernel[7]+tmp[3003]*kernel[8];
				ans[2903]<=tmp[2802]*kernel[0]+tmp[2803]*kernel[1]+tmp[2804]*kernel[2]+tmp[2902]*kernel[3]+tmp[2903]*kernel[4]+tmp[2904]*kernel[5]+tmp[3002]*kernel[6]+tmp[3003]*kernel[7]+tmp[3004]*kernel[8];
				ans[2904]<=tmp[2803]*kernel[0]+tmp[2804]*kernel[1]+tmp[2805]*kernel[2]+tmp[2903]*kernel[3]+tmp[2904]*kernel[4]+tmp[2905]*kernel[5]+tmp[3003]*kernel[6]+tmp[3004]*kernel[7]+tmp[3005]*kernel[8];
				ans[2905]<=tmp[2804]*kernel[0]+tmp[2805]*kernel[1]+tmp[2806]*kernel[2]+tmp[2904]*kernel[3]+tmp[2905]*kernel[4]+tmp[2906]*kernel[5]+tmp[3004]*kernel[6]+tmp[3005]*kernel[7]+tmp[3006]*kernel[8];
				ans[2906]<=tmp[2805]*kernel[0]+tmp[2806]*kernel[1]+tmp[2807]*kernel[2]+tmp[2905]*kernel[3]+tmp[2906]*kernel[4]+tmp[2907]*kernel[5]+tmp[3005]*kernel[6]+tmp[3006]*kernel[7]+tmp[3007]*kernel[8];
				ans[2907]<=tmp[2806]*kernel[0]+tmp[2807]*kernel[1]+tmp[2808]*kernel[2]+tmp[2906]*kernel[3]+tmp[2907]*kernel[4]+tmp[2908]*kernel[5]+tmp[3006]*kernel[6]+tmp[3007]*kernel[7]+tmp[3008]*kernel[8];
				ans[2908]<=tmp[2807]*kernel[0]+tmp[2808]*kernel[1]+tmp[2809]*kernel[2]+tmp[2907]*kernel[3]+tmp[2908]*kernel[4]+tmp[2909]*kernel[5]+tmp[3007]*kernel[6]+tmp[3008]*kernel[7]+tmp[3009]*kernel[8];
				ans[2909]<=tmp[2808]*kernel[0]+tmp[2809]*kernel[1]+tmp[2810]*kernel[2]+tmp[2908]*kernel[3]+tmp[2909]*kernel[4]+tmp[2910]*kernel[5]+tmp[3008]*kernel[6]+tmp[3009]*kernel[7]+tmp[3010]*kernel[8];
				ans[2910]<=tmp[2809]*kernel[0]+tmp[2810]*kernel[1]+tmp[2811]*kernel[2]+tmp[2909]*kernel[3]+tmp[2910]*kernel[4]+tmp[2911]*kernel[5]+tmp[3009]*kernel[6]+tmp[3010]*kernel[7]+tmp[3011]*kernel[8];
				ans[2911]<=tmp[2810]*kernel[0]+tmp[2811]*kernel[1]+tmp[2812]*kernel[2]+tmp[2910]*kernel[3]+tmp[2911]*kernel[4]+tmp[2912]*kernel[5]+tmp[3010]*kernel[6]+tmp[3011]*kernel[7]+tmp[3012]*kernel[8];
				ans[2912]<=tmp[2811]*kernel[0]+tmp[2812]*kernel[1]+tmp[2813]*kernel[2]+tmp[2911]*kernel[3]+tmp[2912]*kernel[4]+tmp[2913]*kernel[5]+tmp[3011]*kernel[6]+tmp[3012]*kernel[7]+tmp[3013]*kernel[8];
				ans[2913]<=tmp[2812]*kernel[0]+tmp[2813]*kernel[1]+tmp[2814]*kernel[2]+tmp[2912]*kernel[3]+tmp[2913]*kernel[4]+tmp[2914]*kernel[5]+tmp[3012]*kernel[6]+tmp[3013]*kernel[7]+tmp[3014]*kernel[8];
				ans[2914]<=tmp[2813]*kernel[0]+tmp[2814]*kernel[1]+tmp[2815]*kernel[2]+tmp[2913]*kernel[3]+tmp[2914]*kernel[4]+tmp[2915]*kernel[5]+tmp[3013]*kernel[6]+tmp[3014]*kernel[7]+tmp[3015]*kernel[8];
				ans[2915]<=tmp[2814]*kernel[0]+tmp[2815]*kernel[1]+tmp[2816]*kernel[2]+tmp[2914]*kernel[3]+tmp[2915]*kernel[4]+tmp[2916]*kernel[5]+tmp[3014]*kernel[6]+tmp[3015]*kernel[7]+tmp[3016]*kernel[8];
				ans[2916]<=tmp[2815]*kernel[0]+tmp[2816]*kernel[1]+tmp[2817]*kernel[2]+tmp[2915]*kernel[3]+tmp[2916]*kernel[4]+tmp[2917]*kernel[5]+tmp[3015]*kernel[6]+tmp[3016]*kernel[7]+tmp[3017]*kernel[8];
				ans[2917]<=tmp[2816]*kernel[0]+tmp[2817]*kernel[1]+tmp[2818]*kernel[2]+tmp[2916]*kernel[3]+tmp[2917]*kernel[4]+tmp[2918]*kernel[5]+tmp[3016]*kernel[6]+tmp[3017]*kernel[7]+tmp[3018]*kernel[8];
				ans[2918]<=tmp[2817]*kernel[0]+tmp[2818]*kernel[1]+tmp[2819]*kernel[2]+tmp[2917]*kernel[3]+tmp[2918]*kernel[4]+tmp[2919]*kernel[5]+tmp[3017]*kernel[6]+tmp[3018]*kernel[7]+tmp[3019]*kernel[8];
				ans[2919]<=tmp[2818]*kernel[0]+tmp[2819]*kernel[1]+tmp[2820]*kernel[2]+tmp[2918]*kernel[3]+tmp[2919]*kernel[4]+tmp[2920]*kernel[5]+tmp[3018]*kernel[6]+tmp[3019]*kernel[7]+tmp[3020]*kernel[8];
				ans[2920]<=tmp[2819]*kernel[0]+tmp[2820]*kernel[1]+tmp[2821]*kernel[2]+tmp[2919]*kernel[3]+tmp[2920]*kernel[4]+tmp[2921]*kernel[5]+tmp[3019]*kernel[6]+tmp[3020]*kernel[7]+tmp[3021]*kernel[8];
				ans[2921]<=tmp[2820]*kernel[0]+tmp[2821]*kernel[1]+tmp[2822]*kernel[2]+tmp[2920]*kernel[3]+tmp[2921]*kernel[4]+tmp[2922]*kernel[5]+tmp[3020]*kernel[6]+tmp[3021]*kernel[7]+tmp[3022]*kernel[8];
				ans[2922]<=tmp[2821]*kernel[0]+tmp[2822]*kernel[1]+tmp[2823]*kernel[2]+tmp[2921]*kernel[3]+tmp[2922]*kernel[4]+tmp[2923]*kernel[5]+tmp[3021]*kernel[6]+tmp[3022]*kernel[7]+tmp[3023]*kernel[8];
				ans[2923]<=tmp[2822]*kernel[0]+tmp[2823]*kernel[1]+tmp[2824]*kernel[2]+tmp[2922]*kernel[3]+tmp[2923]*kernel[4]+tmp[2924]*kernel[5]+tmp[3022]*kernel[6]+tmp[3023]*kernel[7]+tmp[3024]*kernel[8];
				ans[2924]<=tmp[2823]*kernel[0]+tmp[2824]*kernel[1]+tmp[2825]*kernel[2]+tmp[2923]*kernel[3]+tmp[2924]*kernel[4]+tmp[2925]*kernel[5]+tmp[3023]*kernel[6]+tmp[3024]*kernel[7]+tmp[3025]*kernel[8];
				ans[2925]<=tmp[2824]*kernel[0]+tmp[2825]*kernel[1]+tmp[2826]*kernel[2]+tmp[2924]*kernel[3]+tmp[2925]*kernel[4]+tmp[2926]*kernel[5]+tmp[3024]*kernel[6]+tmp[3025]*kernel[7]+tmp[3026]*kernel[8];
				ans[2926]<=tmp[2825]*kernel[0]+tmp[2826]*kernel[1]+tmp[2827]*kernel[2]+tmp[2925]*kernel[3]+tmp[2926]*kernel[4]+tmp[2927]*kernel[5]+tmp[3025]*kernel[6]+tmp[3026]*kernel[7]+tmp[3027]*kernel[8];
				ans[2927]<=tmp[2826]*kernel[0]+tmp[2827]*kernel[1]+tmp[2828]*kernel[2]+tmp[2926]*kernel[3]+tmp[2927]*kernel[4]+tmp[2928]*kernel[5]+tmp[3026]*kernel[6]+tmp[3027]*kernel[7]+tmp[3028]*kernel[8];
				ans[2928]<=tmp[2827]*kernel[0]+tmp[2828]*kernel[1]+tmp[2829]*kernel[2]+tmp[2927]*kernel[3]+tmp[2928]*kernel[4]+tmp[2929]*kernel[5]+tmp[3027]*kernel[6]+tmp[3028]*kernel[7]+tmp[3029]*kernel[8];
				ans[2929]<=tmp[2828]*kernel[0]+tmp[2829]*kernel[1]+tmp[2830]*kernel[2]+tmp[2928]*kernel[3]+tmp[2929]*kernel[4]+tmp[2930]*kernel[5]+tmp[3028]*kernel[6]+tmp[3029]*kernel[7]+tmp[3030]*kernel[8];
				ans[2930]<=tmp[2829]*kernel[0]+tmp[2830]*kernel[1]+tmp[2831]*kernel[2]+tmp[2929]*kernel[3]+tmp[2930]*kernel[4]+tmp[2931]*kernel[5]+tmp[3029]*kernel[6]+tmp[3030]*kernel[7]+tmp[3031]*kernel[8];
				ans[2931]<=tmp[2830]*kernel[0]+tmp[2831]*kernel[1]+tmp[2832]*kernel[2]+tmp[2930]*kernel[3]+tmp[2931]*kernel[4]+tmp[2932]*kernel[5]+tmp[3030]*kernel[6]+tmp[3031]*kernel[7]+tmp[3032]*kernel[8];
				ans[2932]<=tmp[2831]*kernel[0]+tmp[2832]*kernel[1]+tmp[2833]*kernel[2]+tmp[2931]*kernel[3]+tmp[2932]*kernel[4]+tmp[2933]*kernel[5]+tmp[3031]*kernel[6]+tmp[3032]*kernel[7]+tmp[3033]*kernel[8];
				ans[2933]<=tmp[2832]*kernel[0]+tmp[2833]*kernel[1]+tmp[2834]*kernel[2]+tmp[2932]*kernel[3]+tmp[2933]*kernel[4]+tmp[2934]*kernel[5]+tmp[3032]*kernel[6]+tmp[3033]*kernel[7]+tmp[3034]*kernel[8];
				ans[2934]<=tmp[2833]*kernel[0]+tmp[2834]*kernel[1]+tmp[2835]*kernel[2]+tmp[2933]*kernel[3]+tmp[2934]*kernel[4]+tmp[2935]*kernel[5]+tmp[3033]*kernel[6]+tmp[3034]*kernel[7]+tmp[3035]*kernel[8];
				ans[2935]<=tmp[2834]*kernel[0]+tmp[2835]*kernel[1]+tmp[2836]*kernel[2]+tmp[2934]*kernel[3]+tmp[2935]*kernel[4]+tmp[2936]*kernel[5]+tmp[3034]*kernel[6]+tmp[3035]*kernel[7]+tmp[3036]*kernel[8];
				ans[2936]<=tmp[2835]*kernel[0]+tmp[2836]*kernel[1]+tmp[2837]*kernel[2]+tmp[2935]*kernel[3]+tmp[2936]*kernel[4]+tmp[2937]*kernel[5]+tmp[3035]*kernel[6]+tmp[3036]*kernel[7]+tmp[3037]*kernel[8];
				ans[2937]<=tmp[2836]*kernel[0]+tmp[2837]*kernel[1]+tmp[2838]*kernel[2]+tmp[2936]*kernel[3]+tmp[2937]*kernel[4]+tmp[2938]*kernel[5]+tmp[3036]*kernel[6]+tmp[3037]*kernel[7]+tmp[3038]*kernel[8];
				ans[2938]<=tmp[2837]*kernel[0]+tmp[2838]*kernel[1]+tmp[2839]*kernel[2]+tmp[2937]*kernel[3]+tmp[2938]*kernel[4]+tmp[2939]*kernel[5]+tmp[3037]*kernel[6]+tmp[3038]*kernel[7]+tmp[3039]*kernel[8];
				ans[2939]<=tmp[2838]*kernel[0]+tmp[2839]*kernel[1]+tmp[2840]*kernel[2]+tmp[2938]*kernel[3]+tmp[2939]*kernel[4]+tmp[2940]*kernel[5]+tmp[3038]*kernel[6]+tmp[3039]*kernel[7]+tmp[3040]*kernel[8];
				ans[2940]<=tmp[2839]*kernel[0]+tmp[2840]*kernel[1]+tmp[2841]*kernel[2]+tmp[2939]*kernel[3]+tmp[2940]*kernel[4]+tmp[2941]*kernel[5]+tmp[3039]*kernel[6]+tmp[3040]*kernel[7]+tmp[3041]*kernel[8];
				ans[2941]<=tmp[2840]*kernel[0]+tmp[2841]*kernel[1]+tmp[2842]*kernel[2]+tmp[2940]*kernel[3]+tmp[2941]*kernel[4]+tmp[2942]*kernel[5]+tmp[3040]*kernel[6]+tmp[3041]*kernel[7]+tmp[3042]*kernel[8];
				ans[2942]<=tmp[2841]*kernel[0]+tmp[2842]*kernel[1]+tmp[2843]*kernel[2]+tmp[2941]*kernel[3]+tmp[2942]*kernel[4]+tmp[2943]*kernel[5]+tmp[3041]*kernel[6]+tmp[3042]*kernel[7]+tmp[3043]*kernel[8];
				ans[2943]<=tmp[2842]*kernel[0]+tmp[2843]*kernel[1]+tmp[2844]*kernel[2]+tmp[2942]*kernel[3]+tmp[2943]*kernel[4]+tmp[2944]*kernel[5]+tmp[3042]*kernel[6]+tmp[3043]*kernel[7]+tmp[3044]*kernel[8];
				ans[2944]<=tmp[2843]*kernel[0]+tmp[2844]*kernel[1]+tmp[2845]*kernel[2]+tmp[2943]*kernel[3]+tmp[2944]*kernel[4]+tmp[2945]*kernel[5]+tmp[3043]*kernel[6]+tmp[3044]*kernel[7]+tmp[3045]*kernel[8];
				ans[2945]<=tmp[2844]*kernel[0]+tmp[2845]*kernel[1]+tmp[2846]*kernel[2]+tmp[2944]*kernel[3]+tmp[2945]*kernel[4]+tmp[2946]*kernel[5]+tmp[3044]*kernel[6]+tmp[3045]*kernel[7]+tmp[3046]*kernel[8];
				ans[2946]<=tmp[2845]*kernel[0]+tmp[2846]*kernel[1]+tmp[2847]*kernel[2]+tmp[2945]*kernel[3]+tmp[2946]*kernel[4]+tmp[2947]*kernel[5]+tmp[3045]*kernel[6]+tmp[3046]*kernel[7]+tmp[3047]*kernel[8];
				ans[2947]<=tmp[2846]*kernel[0]+tmp[2847]*kernel[1]+tmp[2848]*kernel[2]+tmp[2946]*kernel[3]+tmp[2947]*kernel[4]+tmp[2948]*kernel[5]+tmp[3046]*kernel[6]+tmp[3047]*kernel[7]+tmp[3048]*kernel[8];
				ans[2948]<=tmp[2847]*kernel[0]+tmp[2848]*kernel[1]+tmp[2849]*kernel[2]+tmp[2947]*kernel[3]+tmp[2948]*kernel[4]+tmp[2949]*kernel[5]+tmp[3047]*kernel[6]+tmp[3048]*kernel[7]+tmp[3049]*kernel[8];
				ans[2949]<=tmp[2848]*kernel[0]+tmp[2849]*kernel[1]+tmp[2850]*kernel[2]+tmp[2948]*kernel[3]+tmp[2949]*kernel[4]+tmp[2950]*kernel[5]+tmp[3048]*kernel[6]+tmp[3049]*kernel[7]+tmp[3050]*kernel[8];
				ans[2950]<=tmp[2849]*kernel[0]+tmp[2850]*kernel[1]+tmp[2851]*kernel[2]+tmp[2949]*kernel[3]+tmp[2950]*kernel[4]+tmp[2951]*kernel[5]+tmp[3049]*kernel[6]+tmp[3050]*kernel[7]+tmp[3051]*kernel[8];
				ans[2951]<=tmp[2850]*kernel[0]+tmp[2851]*kernel[1]+tmp[2852]*kernel[2]+tmp[2950]*kernel[3]+tmp[2951]*kernel[4]+tmp[2952]*kernel[5]+tmp[3050]*kernel[6]+tmp[3051]*kernel[7]+tmp[3052]*kernel[8];
				ans[2952]<=tmp[2851]*kernel[0]+tmp[2852]*kernel[1]+tmp[2853]*kernel[2]+tmp[2951]*kernel[3]+tmp[2952]*kernel[4]+tmp[2953]*kernel[5]+tmp[3051]*kernel[6]+tmp[3052]*kernel[7]+tmp[3053]*kernel[8];
				ans[2953]<=tmp[2852]*kernel[0]+tmp[2853]*kernel[1]+tmp[2854]*kernel[2]+tmp[2952]*kernel[3]+tmp[2953]*kernel[4]+tmp[2954]*kernel[5]+tmp[3052]*kernel[6]+tmp[3053]*kernel[7]+tmp[3054]*kernel[8];
				ans[2954]<=tmp[2853]*kernel[0]+tmp[2854]*kernel[1]+tmp[2855]*kernel[2]+tmp[2953]*kernel[3]+tmp[2954]*kernel[4]+tmp[2955]*kernel[5]+tmp[3053]*kernel[6]+tmp[3054]*kernel[7]+tmp[3055]*kernel[8];
				ans[2955]<=tmp[2854]*kernel[0]+tmp[2855]*kernel[1]+tmp[2856]*kernel[2]+tmp[2954]*kernel[3]+tmp[2955]*kernel[4]+tmp[2956]*kernel[5]+tmp[3054]*kernel[6]+tmp[3055]*kernel[7]+tmp[3056]*kernel[8];
				ans[2956]<=tmp[2855]*kernel[0]+tmp[2856]*kernel[1]+tmp[2857]*kernel[2]+tmp[2955]*kernel[3]+tmp[2956]*kernel[4]+tmp[2957]*kernel[5]+tmp[3055]*kernel[6]+tmp[3056]*kernel[7]+tmp[3057]*kernel[8];
				ans[2957]<=tmp[2856]*kernel[0]+tmp[2857]*kernel[1]+tmp[2858]*kernel[2]+tmp[2956]*kernel[3]+tmp[2957]*kernel[4]+tmp[2958]*kernel[5]+tmp[3056]*kernel[6]+tmp[3057]*kernel[7]+tmp[3058]*kernel[8];
				ans[2958]<=tmp[2857]*kernel[0]+tmp[2858]*kernel[1]+tmp[2859]*kernel[2]+tmp[2957]*kernel[3]+tmp[2958]*kernel[4]+tmp[2959]*kernel[5]+tmp[3057]*kernel[6]+tmp[3058]*kernel[7]+tmp[3059]*kernel[8];
				ans[2959]<=tmp[2858]*kernel[0]+tmp[2859]*kernel[1]+tmp[2860]*kernel[2]+tmp[2958]*kernel[3]+tmp[2959]*kernel[4]+tmp[2960]*kernel[5]+tmp[3058]*kernel[6]+tmp[3059]*kernel[7]+tmp[3060]*kernel[8];
				ans[2960]<=tmp[2859]*kernel[0]+tmp[2860]*kernel[1]+tmp[2861]*kernel[2]+tmp[2959]*kernel[3]+tmp[2960]*kernel[4]+tmp[2961]*kernel[5]+tmp[3059]*kernel[6]+tmp[3060]*kernel[7]+tmp[3061]*kernel[8];
				ans[2961]<=tmp[2860]*kernel[0]+tmp[2861]*kernel[1]+tmp[2862]*kernel[2]+tmp[2960]*kernel[3]+tmp[2961]*kernel[4]+tmp[2962]*kernel[5]+tmp[3060]*kernel[6]+tmp[3061]*kernel[7]+tmp[3062]*kernel[8];
				ans[2962]<=tmp[2861]*kernel[0]+tmp[2862]*kernel[1]+tmp[2863]*kernel[2]+tmp[2961]*kernel[3]+tmp[2962]*kernel[4]+tmp[2963]*kernel[5]+tmp[3061]*kernel[6]+tmp[3062]*kernel[7]+tmp[3063]*kernel[8];
				ans[2963]<=tmp[2862]*kernel[0]+tmp[2863]*kernel[1]+tmp[2864]*kernel[2]+tmp[2962]*kernel[3]+tmp[2963]*kernel[4]+tmp[2964]*kernel[5]+tmp[3062]*kernel[6]+tmp[3063]*kernel[7]+tmp[3064]*kernel[8];
				ans[2964]<=tmp[2863]*kernel[0]+tmp[2864]*kernel[1]+tmp[2865]*kernel[2]+tmp[2963]*kernel[3]+tmp[2964]*kernel[4]+tmp[2965]*kernel[5]+tmp[3063]*kernel[6]+tmp[3064]*kernel[7]+tmp[3065]*kernel[8];
				ans[2965]<=tmp[2864]*kernel[0]+tmp[2865]*kernel[1]+tmp[2866]*kernel[2]+tmp[2964]*kernel[3]+tmp[2965]*kernel[4]+tmp[2966]*kernel[5]+tmp[3064]*kernel[6]+tmp[3065]*kernel[7]+tmp[3066]*kernel[8];
				ans[2966]<=tmp[2865]*kernel[0]+tmp[2866]*kernel[1]+tmp[2867]*kernel[2]+tmp[2965]*kernel[3]+tmp[2966]*kernel[4]+tmp[2967]*kernel[5]+tmp[3065]*kernel[6]+tmp[3066]*kernel[7]+tmp[3067]*kernel[8];
				ans[2967]<=tmp[2866]*kernel[0]+tmp[2867]*kernel[1]+tmp[2868]*kernel[2]+tmp[2966]*kernel[3]+tmp[2967]*kernel[4]+tmp[2968]*kernel[5]+tmp[3066]*kernel[6]+tmp[3067]*kernel[7]+tmp[3068]*kernel[8];
				ans[2968]<=tmp[2867]*kernel[0]+tmp[2868]*kernel[1]+tmp[2869]*kernel[2]+tmp[2967]*kernel[3]+tmp[2968]*kernel[4]+tmp[2969]*kernel[5]+tmp[3067]*kernel[6]+tmp[3068]*kernel[7]+tmp[3069]*kernel[8];
				ans[2969]<=tmp[2868]*kernel[0]+tmp[2869]*kernel[1]+tmp[2870]*kernel[2]+tmp[2968]*kernel[3]+tmp[2969]*kernel[4]+tmp[2970]*kernel[5]+tmp[3068]*kernel[6]+tmp[3069]*kernel[7]+tmp[3070]*kernel[8];
				ans[2970]<=tmp[2869]*kernel[0]+tmp[2870]*kernel[1]+tmp[2871]*kernel[2]+tmp[2969]*kernel[3]+tmp[2970]*kernel[4]+tmp[2971]*kernel[5]+tmp[3069]*kernel[6]+tmp[3070]*kernel[7]+tmp[3071]*kernel[8];
				ans[2971]<=tmp[2870]*kernel[0]+tmp[2871]*kernel[1]+tmp[2872]*kernel[2]+tmp[2970]*kernel[3]+tmp[2971]*kernel[4]+tmp[2972]*kernel[5]+tmp[3070]*kernel[6]+tmp[3071]*kernel[7]+tmp[3072]*kernel[8];
				ans[2972]<=tmp[2871]*kernel[0]+tmp[2872]*kernel[1]+tmp[2873]*kernel[2]+tmp[2971]*kernel[3]+tmp[2972]*kernel[4]+tmp[2973]*kernel[5]+tmp[3071]*kernel[6]+tmp[3072]*kernel[7]+tmp[3073]*kernel[8];
				ans[2973]<=tmp[2872]*kernel[0]+tmp[2873]*kernel[1]+tmp[2874]*kernel[2]+tmp[2972]*kernel[3]+tmp[2973]*kernel[4]+tmp[2974]*kernel[5]+tmp[3072]*kernel[6]+tmp[3073]*kernel[7]+tmp[3074]*kernel[8];
				ans[2974]<=tmp[2873]*kernel[0]+tmp[2874]*kernel[1]+tmp[2875]*kernel[2]+tmp[2973]*kernel[3]+tmp[2974]*kernel[4]+tmp[2975]*kernel[5]+tmp[3073]*kernel[6]+tmp[3074]*kernel[7]+tmp[3075]*kernel[8];
				ans[2975]<=tmp[2874]*kernel[0]+tmp[2875]*kernel[1]+tmp[2876]*kernel[2]+tmp[2974]*kernel[3]+tmp[2975]*kernel[4]+tmp[2976]*kernel[5]+tmp[3074]*kernel[6]+tmp[3075]*kernel[7]+tmp[3076]*kernel[8];
				ans[2976]<=tmp[2875]*kernel[0]+tmp[2876]*kernel[1]+tmp[2877]*kernel[2]+tmp[2975]*kernel[3]+tmp[2976]*kernel[4]+tmp[2977]*kernel[5]+tmp[3075]*kernel[6]+tmp[3076]*kernel[7]+tmp[3077]*kernel[8];
				ans[2977]<=tmp[2876]*kernel[0]+tmp[2877]*kernel[1]+tmp[2878]*kernel[2]+tmp[2976]*kernel[3]+tmp[2977]*kernel[4]+tmp[2978]*kernel[5]+tmp[3076]*kernel[6]+tmp[3077]*kernel[7]+tmp[3078]*kernel[8];
				ans[2978]<=tmp[2877]*kernel[0]+tmp[2878]*kernel[1]+tmp[2879]*kernel[2]+tmp[2977]*kernel[3]+tmp[2978]*kernel[4]+tmp[2979]*kernel[5]+tmp[3077]*kernel[6]+tmp[3078]*kernel[7]+tmp[3079]*kernel[8];
				ans[2979]<=tmp[2878]*kernel[0]+tmp[2879]*kernel[1]+tmp[2880]*kernel[2]+tmp[2978]*kernel[3]+tmp[2979]*kernel[4]+tmp[2980]*kernel[5]+tmp[3078]*kernel[6]+tmp[3079]*kernel[7]+tmp[3080]*kernel[8];
				ans[2980]<=tmp[2879]*kernel[0]+tmp[2880]*kernel[1]+tmp[2881]*kernel[2]+tmp[2979]*kernel[3]+tmp[2980]*kernel[4]+tmp[2981]*kernel[5]+tmp[3079]*kernel[6]+tmp[3080]*kernel[7]+tmp[3081]*kernel[8];
				ans[2981]<=tmp[2880]*kernel[0]+tmp[2881]*kernel[1]+tmp[2882]*kernel[2]+tmp[2980]*kernel[3]+tmp[2981]*kernel[4]+tmp[2982]*kernel[5]+tmp[3080]*kernel[6]+tmp[3081]*kernel[7]+tmp[3082]*kernel[8];
				ans[2982]<=tmp[2881]*kernel[0]+tmp[2882]*kernel[1]+tmp[2883]*kernel[2]+tmp[2981]*kernel[3]+tmp[2982]*kernel[4]+tmp[2983]*kernel[5]+tmp[3081]*kernel[6]+tmp[3082]*kernel[7]+tmp[3083]*kernel[8];
				ans[2983]<=tmp[2882]*kernel[0]+tmp[2883]*kernel[1]+tmp[2884]*kernel[2]+tmp[2982]*kernel[3]+tmp[2983]*kernel[4]+tmp[2984]*kernel[5]+tmp[3082]*kernel[6]+tmp[3083]*kernel[7]+tmp[3084]*kernel[8];
				ans[2984]<=tmp[2883]*kernel[0]+tmp[2884]*kernel[1]+tmp[2885]*kernel[2]+tmp[2983]*kernel[3]+tmp[2984]*kernel[4]+tmp[2985]*kernel[5]+tmp[3083]*kernel[6]+tmp[3084]*kernel[7]+tmp[3085]*kernel[8];
				ans[2985]<=tmp[2884]*kernel[0]+tmp[2885]*kernel[1]+tmp[2886]*kernel[2]+tmp[2984]*kernel[3]+tmp[2985]*kernel[4]+tmp[2986]*kernel[5]+tmp[3084]*kernel[6]+tmp[3085]*kernel[7]+tmp[3086]*kernel[8];
				ans[2986]<=tmp[2885]*kernel[0]+tmp[2886]*kernel[1]+tmp[2887]*kernel[2]+tmp[2985]*kernel[3]+tmp[2986]*kernel[4]+tmp[2987]*kernel[5]+tmp[3085]*kernel[6]+tmp[3086]*kernel[7]+tmp[3087]*kernel[8];
				ans[2987]<=tmp[2886]*kernel[0]+tmp[2887]*kernel[1]+tmp[2888]*kernel[2]+tmp[2986]*kernel[3]+tmp[2987]*kernel[4]+tmp[2988]*kernel[5]+tmp[3086]*kernel[6]+tmp[3087]*kernel[7]+tmp[3088]*kernel[8];
				ans[2988]<=tmp[2887]*kernel[0]+tmp[2888]*kernel[1]+tmp[2889]*kernel[2]+tmp[2987]*kernel[3]+tmp[2988]*kernel[4]+tmp[2989]*kernel[5]+tmp[3087]*kernel[6]+tmp[3088]*kernel[7]+tmp[3089]*kernel[8];
				ans[2989]<=tmp[2888]*kernel[0]+tmp[2889]*kernel[1]+tmp[2890]*kernel[2]+tmp[2988]*kernel[3]+tmp[2989]*kernel[4]+tmp[2990]*kernel[5]+tmp[3088]*kernel[6]+tmp[3089]*kernel[7]+tmp[3090]*kernel[8];
				ans[2990]<=tmp[2889]*kernel[0]+tmp[2890]*kernel[1]+tmp[2891]*kernel[2]+tmp[2989]*kernel[3]+tmp[2990]*kernel[4]+tmp[2991]*kernel[5]+tmp[3089]*kernel[6]+tmp[3090]*kernel[7]+tmp[3091]*kernel[8];
				ans[2991]<=tmp[2890]*kernel[0]+tmp[2891]*kernel[1]+tmp[2892]*kernel[2]+tmp[2990]*kernel[3]+tmp[2991]*kernel[4]+tmp[2992]*kernel[5]+tmp[3090]*kernel[6]+tmp[3091]*kernel[7]+tmp[3092]*kernel[8];
				ans[2992]<=tmp[2891]*kernel[0]+tmp[2892]*kernel[1]+tmp[2893]*kernel[2]+tmp[2991]*kernel[3]+tmp[2992]*kernel[4]+tmp[2993]*kernel[5]+tmp[3091]*kernel[6]+tmp[3092]*kernel[7]+tmp[3093]*kernel[8];
				ans[2993]<=tmp[2892]*kernel[0]+tmp[2893]*kernel[1]+tmp[2894]*kernel[2]+tmp[2992]*kernel[3]+tmp[2993]*kernel[4]+tmp[2994]*kernel[5]+tmp[3092]*kernel[6]+tmp[3093]*kernel[7]+tmp[3094]*kernel[8];
				ans[2994]<=tmp[2893]*kernel[0]+tmp[2894]*kernel[1]+tmp[2895]*kernel[2]+tmp[2993]*kernel[3]+tmp[2994]*kernel[4]+tmp[2995]*kernel[5]+tmp[3093]*kernel[6]+tmp[3094]*kernel[7]+tmp[3095]*kernel[8];
				ans[2995]<=tmp[2894]*kernel[0]+tmp[2895]*kernel[1]+tmp[2896]*kernel[2]+tmp[2994]*kernel[3]+tmp[2995]*kernel[4]+tmp[2996]*kernel[5]+tmp[3094]*kernel[6]+tmp[3095]*kernel[7]+tmp[3096]*kernel[8];
				ans[2996]<=tmp[2895]*kernel[0]+tmp[2896]*kernel[1]+tmp[2897]*kernel[2]+tmp[2995]*kernel[3]+tmp[2996]*kernel[4]+tmp[2997]*kernel[5]+tmp[3095]*kernel[6]+tmp[3096]*kernel[7]+tmp[3097]*kernel[8];
				ans[2997]<=tmp[2896]*kernel[0]+tmp[2897]*kernel[1]+tmp[2898]*kernel[2]+tmp[2996]*kernel[3]+tmp[2997]*kernel[4]+tmp[2998]*kernel[5]+tmp[3096]*kernel[6]+tmp[3097]*kernel[7]+tmp[3098]*kernel[8];
				ans[2998]<=tmp[2897]*kernel[0]+tmp[2898]*kernel[1]+tmp[2899]*kernel[2]+tmp[2997]*kernel[3]+tmp[2998]*kernel[4]+tmp[2999]*kernel[5]+tmp[3097]*kernel[6]+tmp[3098]*kernel[7]+tmp[3099]*kernel[8];
				ans[2999]<=tmp[2898]*kernel[0]+tmp[2899]*kernel[1]+tmp[2998]*kernel[3]+tmp[2999]*kernel[4]+tmp[3098]*kernel[6]+tmp[3099]*kernel[7];
				ans[3000]<=tmp[2900]*kernel[1]+tmp[2901]*kernel[2]+tmp[3000]*kernel[4]+tmp[3001]*kernel[5]+tmp[3100]*kernel[7]+tmp[3101]*kernel[8];
				ans[3001]<=tmp[2900]*kernel[0]+tmp[2901]*kernel[1]+tmp[2902]*kernel[2]+tmp[3000]*kernel[3]+tmp[3001]*kernel[4]+tmp[3002]*kernel[5]+tmp[3100]*kernel[6]+tmp[3101]*kernel[7]+tmp[3102]*kernel[8];
				ans[3002]<=tmp[2901]*kernel[0]+tmp[2902]*kernel[1]+tmp[2903]*kernel[2]+tmp[3001]*kernel[3]+tmp[3002]*kernel[4]+tmp[3003]*kernel[5]+tmp[3101]*kernel[6]+tmp[3102]*kernel[7]+tmp[3103]*kernel[8];
				ans[3003]<=tmp[2902]*kernel[0]+tmp[2903]*kernel[1]+tmp[2904]*kernel[2]+tmp[3002]*kernel[3]+tmp[3003]*kernel[4]+tmp[3004]*kernel[5]+tmp[3102]*kernel[6]+tmp[3103]*kernel[7]+tmp[3104]*kernel[8];
				ans[3004]<=tmp[2903]*kernel[0]+tmp[2904]*kernel[1]+tmp[2905]*kernel[2]+tmp[3003]*kernel[3]+tmp[3004]*kernel[4]+tmp[3005]*kernel[5]+tmp[3103]*kernel[6]+tmp[3104]*kernel[7]+tmp[3105]*kernel[8];
				ans[3005]<=tmp[2904]*kernel[0]+tmp[2905]*kernel[1]+tmp[2906]*kernel[2]+tmp[3004]*kernel[3]+tmp[3005]*kernel[4]+tmp[3006]*kernel[5]+tmp[3104]*kernel[6]+tmp[3105]*kernel[7]+tmp[3106]*kernel[8];
				ans[3006]<=tmp[2905]*kernel[0]+tmp[2906]*kernel[1]+tmp[2907]*kernel[2]+tmp[3005]*kernel[3]+tmp[3006]*kernel[4]+tmp[3007]*kernel[5]+tmp[3105]*kernel[6]+tmp[3106]*kernel[7]+tmp[3107]*kernel[8];
				ans[3007]<=tmp[2906]*kernel[0]+tmp[2907]*kernel[1]+tmp[2908]*kernel[2]+tmp[3006]*kernel[3]+tmp[3007]*kernel[4]+tmp[3008]*kernel[5]+tmp[3106]*kernel[6]+tmp[3107]*kernel[7]+tmp[3108]*kernel[8];
				ans[3008]<=tmp[2907]*kernel[0]+tmp[2908]*kernel[1]+tmp[2909]*kernel[2]+tmp[3007]*kernel[3]+tmp[3008]*kernel[4]+tmp[3009]*kernel[5]+tmp[3107]*kernel[6]+tmp[3108]*kernel[7]+tmp[3109]*kernel[8];
				ans[3009]<=tmp[2908]*kernel[0]+tmp[2909]*kernel[1]+tmp[2910]*kernel[2]+tmp[3008]*kernel[3]+tmp[3009]*kernel[4]+tmp[3010]*kernel[5]+tmp[3108]*kernel[6]+tmp[3109]*kernel[7]+tmp[3110]*kernel[8];
				ans[3010]<=tmp[2909]*kernel[0]+tmp[2910]*kernel[1]+tmp[2911]*kernel[2]+tmp[3009]*kernel[3]+tmp[3010]*kernel[4]+tmp[3011]*kernel[5]+tmp[3109]*kernel[6]+tmp[3110]*kernel[7]+tmp[3111]*kernel[8];
				ans[3011]<=tmp[2910]*kernel[0]+tmp[2911]*kernel[1]+tmp[2912]*kernel[2]+tmp[3010]*kernel[3]+tmp[3011]*kernel[4]+tmp[3012]*kernel[5]+tmp[3110]*kernel[6]+tmp[3111]*kernel[7]+tmp[3112]*kernel[8];
				ans[3012]<=tmp[2911]*kernel[0]+tmp[2912]*kernel[1]+tmp[2913]*kernel[2]+tmp[3011]*kernel[3]+tmp[3012]*kernel[4]+tmp[3013]*kernel[5]+tmp[3111]*kernel[6]+tmp[3112]*kernel[7]+tmp[3113]*kernel[8];
				ans[3013]<=tmp[2912]*kernel[0]+tmp[2913]*kernel[1]+tmp[2914]*kernel[2]+tmp[3012]*kernel[3]+tmp[3013]*kernel[4]+tmp[3014]*kernel[5]+tmp[3112]*kernel[6]+tmp[3113]*kernel[7]+tmp[3114]*kernel[8];
				ans[3014]<=tmp[2913]*kernel[0]+tmp[2914]*kernel[1]+tmp[2915]*kernel[2]+tmp[3013]*kernel[3]+tmp[3014]*kernel[4]+tmp[3015]*kernel[5]+tmp[3113]*kernel[6]+tmp[3114]*kernel[7]+tmp[3115]*kernel[8];
				ans[3015]<=tmp[2914]*kernel[0]+tmp[2915]*kernel[1]+tmp[2916]*kernel[2]+tmp[3014]*kernel[3]+tmp[3015]*kernel[4]+tmp[3016]*kernel[5]+tmp[3114]*kernel[6]+tmp[3115]*kernel[7]+tmp[3116]*kernel[8];
				ans[3016]<=tmp[2915]*kernel[0]+tmp[2916]*kernel[1]+tmp[2917]*kernel[2]+tmp[3015]*kernel[3]+tmp[3016]*kernel[4]+tmp[3017]*kernel[5]+tmp[3115]*kernel[6]+tmp[3116]*kernel[7]+tmp[3117]*kernel[8];
				ans[3017]<=tmp[2916]*kernel[0]+tmp[2917]*kernel[1]+tmp[2918]*kernel[2]+tmp[3016]*kernel[3]+tmp[3017]*kernel[4]+tmp[3018]*kernel[5]+tmp[3116]*kernel[6]+tmp[3117]*kernel[7]+tmp[3118]*kernel[8];
				ans[3018]<=tmp[2917]*kernel[0]+tmp[2918]*kernel[1]+tmp[2919]*kernel[2]+tmp[3017]*kernel[3]+tmp[3018]*kernel[4]+tmp[3019]*kernel[5]+tmp[3117]*kernel[6]+tmp[3118]*kernel[7]+tmp[3119]*kernel[8];
				ans[3019]<=tmp[2918]*kernel[0]+tmp[2919]*kernel[1]+tmp[2920]*kernel[2]+tmp[3018]*kernel[3]+tmp[3019]*kernel[4]+tmp[3020]*kernel[5]+tmp[3118]*kernel[6]+tmp[3119]*kernel[7]+tmp[3120]*kernel[8];
				ans[3020]<=tmp[2919]*kernel[0]+tmp[2920]*kernel[1]+tmp[2921]*kernel[2]+tmp[3019]*kernel[3]+tmp[3020]*kernel[4]+tmp[3021]*kernel[5]+tmp[3119]*kernel[6]+tmp[3120]*kernel[7]+tmp[3121]*kernel[8];
				ans[3021]<=tmp[2920]*kernel[0]+tmp[2921]*kernel[1]+tmp[2922]*kernel[2]+tmp[3020]*kernel[3]+tmp[3021]*kernel[4]+tmp[3022]*kernel[5]+tmp[3120]*kernel[6]+tmp[3121]*kernel[7]+tmp[3122]*kernel[8];
				ans[3022]<=tmp[2921]*kernel[0]+tmp[2922]*kernel[1]+tmp[2923]*kernel[2]+tmp[3021]*kernel[3]+tmp[3022]*kernel[4]+tmp[3023]*kernel[5]+tmp[3121]*kernel[6]+tmp[3122]*kernel[7]+tmp[3123]*kernel[8];
				ans[3023]<=tmp[2922]*kernel[0]+tmp[2923]*kernel[1]+tmp[2924]*kernel[2]+tmp[3022]*kernel[3]+tmp[3023]*kernel[4]+tmp[3024]*kernel[5]+tmp[3122]*kernel[6]+tmp[3123]*kernel[7]+tmp[3124]*kernel[8];
				ans[3024]<=tmp[2923]*kernel[0]+tmp[2924]*kernel[1]+tmp[2925]*kernel[2]+tmp[3023]*kernel[3]+tmp[3024]*kernel[4]+tmp[3025]*kernel[5]+tmp[3123]*kernel[6]+tmp[3124]*kernel[7]+tmp[3125]*kernel[8];
				ans[3025]<=tmp[2924]*kernel[0]+tmp[2925]*kernel[1]+tmp[2926]*kernel[2]+tmp[3024]*kernel[3]+tmp[3025]*kernel[4]+tmp[3026]*kernel[5]+tmp[3124]*kernel[6]+tmp[3125]*kernel[7]+tmp[3126]*kernel[8];
				ans[3026]<=tmp[2925]*kernel[0]+tmp[2926]*kernel[1]+tmp[2927]*kernel[2]+tmp[3025]*kernel[3]+tmp[3026]*kernel[4]+tmp[3027]*kernel[5]+tmp[3125]*kernel[6]+tmp[3126]*kernel[7]+tmp[3127]*kernel[8];
				ans[3027]<=tmp[2926]*kernel[0]+tmp[2927]*kernel[1]+tmp[2928]*kernel[2]+tmp[3026]*kernel[3]+tmp[3027]*kernel[4]+tmp[3028]*kernel[5]+tmp[3126]*kernel[6]+tmp[3127]*kernel[7]+tmp[3128]*kernel[8];
				ans[3028]<=tmp[2927]*kernel[0]+tmp[2928]*kernel[1]+tmp[2929]*kernel[2]+tmp[3027]*kernel[3]+tmp[3028]*kernel[4]+tmp[3029]*kernel[5]+tmp[3127]*kernel[6]+tmp[3128]*kernel[7]+tmp[3129]*kernel[8];
				ans[3029]<=tmp[2928]*kernel[0]+tmp[2929]*kernel[1]+tmp[2930]*kernel[2]+tmp[3028]*kernel[3]+tmp[3029]*kernel[4]+tmp[3030]*kernel[5]+tmp[3128]*kernel[6]+tmp[3129]*kernel[7]+tmp[3130]*kernel[8];
				ans[3030]<=tmp[2929]*kernel[0]+tmp[2930]*kernel[1]+tmp[2931]*kernel[2]+tmp[3029]*kernel[3]+tmp[3030]*kernel[4]+tmp[3031]*kernel[5]+tmp[3129]*kernel[6]+tmp[3130]*kernel[7]+tmp[3131]*kernel[8];
				ans[3031]<=tmp[2930]*kernel[0]+tmp[2931]*kernel[1]+tmp[2932]*kernel[2]+tmp[3030]*kernel[3]+tmp[3031]*kernel[4]+tmp[3032]*kernel[5]+tmp[3130]*kernel[6]+tmp[3131]*kernel[7]+tmp[3132]*kernel[8];
				ans[3032]<=tmp[2931]*kernel[0]+tmp[2932]*kernel[1]+tmp[2933]*kernel[2]+tmp[3031]*kernel[3]+tmp[3032]*kernel[4]+tmp[3033]*kernel[5]+tmp[3131]*kernel[6]+tmp[3132]*kernel[7]+tmp[3133]*kernel[8];
				ans[3033]<=tmp[2932]*kernel[0]+tmp[2933]*kernel[1]+tmp[2934]*kernel[2]+tmp[3032]*kernel[3]+tmp[3033]*kernel[4]+tmp[3034]*kernel[5]+tmp[3132]*kernel[6]+tmp[3133]*kernel[7]+tmp[3134]*kernel[8];
				ans[3034]<=tmp[2933]*kernel[0]+tmp[2934]*kernel[1]+tmp[2935]*kernel[2]+tmp[3033]*kernel[3]+tmp[3034]*kernel[4]+tmp[3035]*kernel[5]+tmp[3133]*kernel[6]+tmp[3134]*kernel[7]+tmp[3135]*kernel[8];
				ans[3035]<=tmp[2934]*kernel[0]+tmp[2935]*kernel[1]+tmp[2936]*kernel[2]+tmp[3034]*kernel[3]+tmp[3035]*kernel[4]+tmp[3036]*kernel[5]+tmp[3134]*kernel[6]+tmp[3135]*kernel[7]+tmp[3136]*kernel[8];
				ans[3036]<=tmp[2935]*kernel[0]+tmp[2936]*kernel[1]+tmp[2937]*kernel[2]+tmp[3035]*kernel[3]+tmp[3036]*kernel[4]+tmp[3037]*kernel[5]+tmp[3135]*kernel[6]+tmp[3136]*kernel[7]+tmp[3137]*kernel[8];
				ans[3037]<=tmp[2936]*kernel[0]+tmp[2937]*kernel[1]+tmp[2938]*kernel[2]+tmp[3036]*kernel[3]+tmp[3037]*kernel[4]+tmp[3038]*kernel[5]+tmp[3136]*kernel[6]+tmp[3137]*kernel[7]+tmp[3138]*kernel[8];
				ans[3038]<=tmp[2937]*kernel[0]+tmp[2938]*kernel[1]+tmp[2939]*kernel[2]+tmp[3037]*kernel[3]+tmp[3038]*kernel[4]+tmp[3039]*kernel[5]+tmp[3137]*kernel[6]+tmp[3138]*kernel[7]+tmp[3139]*kernel[8];
				ans[3039]<=tmp[2938]*kernel[0]+tmp[2939]*kernel[1]+tmp[2940]*kernel[2]+tmp[3038]*kernel[3]+tmp[3039]*kernel[4]+tmp[3040]*kernel[5]+tmp[3138]*kernel[6]+tmp[3139]*kernel[7]+tmp[3140]*kernel[8];
				ans[3040]<=tmp[2939]*kernel[0]+tmp[2940]*kernel[1]+tmp[2941]*kernel[2]+tmp[3039]*kernel[3]+tmp[3040]*kernel[4]+tmp[3041]*kernel[5]+tmp[3139]*kernel[6]+tmp[3140]*kernel[7]+tmp[3141]*kernel[8];
				ans[3041]<=tmp[2940]*kernel[0]+tmp[2941]*kernel[1]+tmp[2942]*kernel[2]+tmp[3040]*kernel[3]+tmp[3041]*kernel[4]+tmp[3042]*kernel[5]+tmp[3140]*kernel[6]+tmp[3141]*kernel[7]+tmp[3142]*kernel[8];
				ans[3042]<=tmp[2941]*kernel[0]+tmp[2942]*kernel[1]+tmp[2943]*kernel[2]+tmp[3041]*kernel[3]+tmp[3042]*kernel[4]+tmp[3043]*kernel[5]+tmp[3141]*kernel[6]+tmp[3142]*kernel[7]+tmp[3143]*kernel[8];
				ans[3043]<=tmp[2942]*kernel[0]+tmp[2943]*kernel[1]+tmp[2944]*kernel[2]+tmp[3042]*kernel[3]+tmp[3043]*kernel[4]+tmp[3044]*kernel[5]+tmp[3142]*kernel[6]+tmp[3143]*kernel[7]+tmp[3144]*kernel[8];
				ans[3044]<=tmp[2943]*kernel[0]+tmp[2944]*kernel[1]+tmp[2945]*kernel[2]+tmp[3043]*kernel[3]+tmp[3044]*kernel[4]+tmp[3045]*kernel[5]+tmp[3143]*kernel[6]+tmp[3144]*kernel[7]+tmp[3145]*kernel[8];
				ans[3045]<=tmp[2944]*kernel[0]+tmp[2945]*kernel[1]+tmp[2946]*kernel[2]+tmp[3044]*kernel[3]+tmp[3045]*kernel[4]+tmp[3046]*kernel[5]+tmp[3144]*kernel[6]+tmp[3145]*kernel[7]+tmp[3146]*kernel[8];
				ans[3046]<=tmp[2945]*kernel[0]+tmp[2946]*kernel[1]+tmp[2947]*kernel[2]+tmp[3045]*kernel[3]+tmp[3046]*kernel[4]+tmp[3047]*kernel[5]+tmp[3145]*kernel[6]+tmp[3146]*kernel[7]+tmp[3147]*kernel[8];
				ans[3047]<=tmp[2946]*kernel[0]+tmp[2947]*kernel[1]+tmp[2948]*kernel[2]+tmp[3046]*kernel[3]+tmp[3047]*kernel[4]+tmp[3048]*kernel[5]+tmp[3146]*kernel[6]+tmp[3147]*kernel[7]+tmp[3148]*kernel[8];
				ans[3048]<=tmp[2947]*kernel[0]+tmp[2948]*kernel[1]+tmp[2949]*kernel[2]+tmp[3047]*kernel[3]+tmp[3048]*kernel[4]+tmp[3049]*kernel[5]+tmp[3147]*kernel[6]+tmp[3148]*kernel[7]+tmp[3149]*kernel[8];
				ans[3049]<=tmp[2948]*kernel[0]+tmp[2949]*kernel[1]+tmp[2950]*kernel[2]+tmp[3048]*kernel[3]+tmp[3049]*kernel[4]+tmp[3050]*kernel[5]+tmp[3148]*kernel[6]+tmp[3149]*kernel[7]+tmp[3150]*kernel[8];
				ans[3050]<=tmp[2949]*kernel[0]+tmp[2950]*kernel[1]+tmp[2951]*kernel[2]+tmp[3049]*kernel[3]+tmp[3050]*kernel[4]+tmp[3051]*kernel[5]+tmp[3149]*kernel[6]+tmp[3150]*kernel[7]+tmp[3151]*kernel[8];
				ans[3051]<=tmp[2950]*kernel[0]+tmp[2951]*kernel[1]+tmp[2952]*kernel[2]+tmp[3050]*kernel[3]+tmp[3051]*kernel[4]+tmp[3052]*kernel[5]+tmp[3150]*kernel[6]+tmp[3151]*kernel[7]+tmp[3152]*kernel[8];
				ans[3052]<=tmp[2951]*kernel[0]+tmp[2952]*kernel[1]+tmp[2953]*kernel[2]+tmp[3051]*kernel[3]+tmp[3052]*kernel[4]+tmp[3053]*kernel[5]+tmp[3151]*kernel[6]+tmp[3152]*kernel[7]+tmp[3153]*kernel[8];
				ans[3053]<=tmp[2952]*kernel[0]+tmp[2953]*kernel[1]+tmp[2954]*kernel[2]+tmp[3052]*kernel[3]+tmp[3053]*kernel[4]+tmp[3054]*kernel[5]+tmp[3152]*kernel[6]+tmp[3153]*kernel[7]+tmp[3154]*kernel[8];
				ans[3054]<=tmp[2953]*kernel[0]+tmp[2954]*kernel[1]+tmp[2955]*kernel[2]+tmp[3053]*kernel[3]+tmp[3054]*kernel[4]+tmp[3055]*kernel[5]+tmp[3153]*kernel[6]+tmp[3154]*kernel[7]+tmp[3155]*kernel[8];
				ans[3055]<=tmp[2954]*kernel[0]+tmp[2955]*kernel[1]+tmp[2956]*kernel[2]+tmp[3054]*kernel[3]+tmp[3055]*kernel[4]+tmp[3056]*kernel[5]+tmp[3154]*kernel[6]+tmp[3155]*kernel[7]+tmp[3156]*kernel[8];
				ans[3056]<=tmp[2955]*kernel[0]+tmp[2956]*kernel[1]+tmp[2957]*kernel[2]+tmp[3055]*kernel[3]+tmp[3056]*kernel[4]+tmp[3057]*kernel[5]+tmp[3155]*kernel[6]+tmp[3156]*kernel[7]+tmp[3157]*kernel[8];
				ans[3057]<=tmp[2956]*kernel[0]+tmp[2957]*kernel[1]+tmp[2958]*kernel[2]+tmp[3056]*kernel[3]+tmp[3057]*kernel[4]+tmp[3058]*kernel[5]+tmp[3156]*kernel[6]+tmp[3157]*kernel[7]+tmp[3158]*kernel[8];
				ans[3058]<=tmp[2957]*kernel[0]+tmp[2958]*kernel[1]+tmp[2959]*kernel[2]+tmp[3057]*kernel[3]+tmp[3058]*kernel[4]+tmp[3059]*kernel[5]+tmp[3157]*kernel[6]+tmp[3158]*kernel[7]+tmp[3159]*kernel[8];
				ans[3059]<=tmp[2958]*kernel[0]+tmp[2959]*kernel[1]+tmp[2960]*kernel[2]+tmp[3058]*kernel[3]+tmp[3059]*kernel[4]+tmp[3060]*kernel[5]+tmp[3158]*kernel[6]+tmp[3159]*kernel[7]+tmp[3160]*kernel[8];
				ans[3060]<=tmp[2959]*kernel[0]+tmp[2960]*kernel[1]+tmp[2961]*kernel[2]+tmp[3059]*kernel[3]+tmp[3060]*kernel[4]+tmp[3061]*kernel[5]+tmp[3159]*kernel[6]+tmp[3160]*kernel[7]+tmp[3161]*kernel[8];
				ans[3061]<=tmp[2960]*kernel[0]+tmp[2961]*kernel[1]+tmp[2962]*kernel[2]+tmp[3060]*kernel[3]+tmp[3061]*kernel[4]+tmp[3062]*kernel[5]+tmp[3160]*kernel[6]+tmp[3161]*kernel[7]+tmp[3162]*kernel[8];
				ans[3062]<=tmp[2961]*kernel[0]+tmp[2962]*kernel[1]+tmp[2963]*kernel[2]+tmp[3061]*kernel[3]+tmp[3062]*kernel[4]+tmp[3063]*kernel[5]+tmp[3161]*kernel[6]+tmp[3162]*kernel[7]+tmp[3163]*kernel[8];
				ans[3063]<=tmp[2962]*kernel[0]+tmp[2963]*kernel[1]+tmp[2964]*kernel[2]+tmp[3062]*kernel[3]+tmp[3063]*kernel[4]+tmp[3064]*kernel[5]+tmp[3162]*kernel[6]+tmp[3163]*kernel[7]+tmp[3164]*kernel[8];
				ans[3064]<=tmp[2963]*kernel[0]+tmp[2964]*kernel[1]+tmp[2965]*kernel[2]+tmp[3063]*kernel[3]+tmp[3064]*kernel[4]+tmp[3065]*kernel[5]+tmp[3163]*kernel[6]+tmp[3164]*kernel[7]+tmp[3165]*kernel[8];
				ans[3065]<=tmp[2964]*kernel[0]+tmp[2965]*kernel[1]+tmp[2966]*kernel[2]+tmp[3064]*kernel[3]+tmp[3065]*kernel[4]+tmp[3066]*kernel[5]+tmp[3164]*kernel[6]+tmp[3165]*kernel[7]+tmp[3166]*kernel[8];
				ans[3066]<=tmp[2965]*kernel[0]+tmp[2966]*kernel[1]+tmp[2967]*kernel[2]+tmp[3065]*kernel[3]+tmp[3066]*kernel[4]+tmp[3067]*kernel[5]+tmp[3165]*kernel[6]+tmp[3166]*kernel[7]+tmp[3167]*kernel[8];
				ans[3067]<=tmp[2966]*kernel[0]+tmp[2967]*kernel[1]+tmp[2968]*kernel[2]+tmp[3066]*kernel[3]+tmp[3067]*kernel[4]+tmp[3068]*kernel[5]+tmp[3166]*kernel[6]+tmp[3167]*kernel[7]+tmp[3168]*kernel[8];
				ans[3068]<=tmp[2967]*kernel[0]+tmp[2968]*kernel[1]+tmp[2969]*kernel[2]+tmp[3067]*kernel[3]+tmp[3068]*kernel[4]+tmp[3069]*kernel[5]+tmp[3167]*kernel[6]+tmp[3168]*kernel[7]+tmp[3169]*kernel[8];
				ans[3069]<=tmp[2968]*kernel[0]+tmp[2969]*kernel[1]+tmp[2970]*kernel[2]+tmp[3068]*kernel[3]+tmp[3069]*kernel[4]+tmp[3070]*kernel[5]+tmp[3168]*kernel[6]+tmp[3169]*kernel[7]+tmp[3170]*kernel[8];
				ans[3070]<=tmp[2969]*kernel[0]+tmp[2970]*kernel[1]+tmp[2971]*kernel[2]+tmp[3069]*kernel[3]+tmp[3070]*kernel[4]+tmp[3071]*kernel[5]+tmp[3169]*kernel[6]+tmp[3170]*kernel[7]+tmp[3171]*kernel[8];
				ans[3071]<=tmp[2970]*kernel[0]+tmp[2971]*kernel[1]+tmp[2972]*kernel[2]+tmp[3070]*kernel[3]+tmp[3071]*kernel[4]+tmp[3072]*kernel[5]+tmp[3170]*kernel[6]+tmp[3171]*kernel[7]+tmp[3172]*kernel[8];
				ans[3072]<=tmp[2971]*kernel[0]+tmp[2972]*kernel[1]+tmp[2973]*kernel[2]+tmp[3071]*kernel[3]+tmp[3072]*kernel[4]+tmp[3073]*kernel[5]+tmp[3171]*kernel[6]+tmp[3172]*kernel[7]+tmp[3173]*kernel[8];
				ans[3073]<=tmp[2972]*kernel[0]+tmp[2973]*kernel[1]+tmp[2974]*kernel[2]+tmp[3072]*kernel[3]+tmp[3073]*kernel[4]+tmp[3074]*kernel[5]+tmp[3172]*kernel[6]+tmp[3173]*kernel[7]+tmp[3174]*kernel[8];
				ans[3074]<=tmp[2973]*kernel[0]+tmp[2974]*kernel[1]+tmp[2975]*kernel[2]+tmp[3073]*kernel[3]+tmp[3074]*kernel[4]+tmp[3075]*kernel[5]+tmp[3173]*kernel[6]+tmp[3174]*kernel[7]+tmp[3175]*kernel[8];
				ans[3075]<=tmp[2974]*kernel[0]+tmp[2975]*kernel[1]+tmp[2976]*kernel[2]+tmp[3074]*kernel[3]+tmp[3075]*kernel[4]+tmp[3076]*kernel[5]+tmp[3174]*kernel[6]+tmp[3175]*kernel[7]+tmp[3176]*kernel[8];
				ans[3076]<=tmp[2975]*kernel[0]+tmp[2976]*kernel[1]+tmp[2977]*kernel[2]+tmp[3075]*kernel[3]+tmp[3076]*kernel[4]+tmp[3077]*kernel[5]+tmp[3175]*kernel[6]+tmp[3176]*kernel[7]+tmp[3177]*kernel[8];
				ans[3077]<=tmp[2976]*kernel[0]+tmp[2977]*kernel[1]+tmp[2978]*kernel[2]+tmp[3076]*kernel[3]+tmp[3077]*kernel[4]+tmp[3078]*kernel[5]+tmp[3176]*kernel[6]+tmp[3177]*kernel[7]+tmp[3178]*kernel[8];
				ans[3078]<=tmp[2977]*kernel[0]+tmp[2978]*kernel[1]+tmp[2979]*kernel[2]+tmp[3077]*kernel[3]+tmp[3078]*kernel[4]+tmp[3079]*kernel[5]+tmp[3177]*kernel[6]+tmp[3178]*kernel[7]+tmp[3179]*kernel[8];
				ans[3079]<=tmp[2978]*kernel[0]+tmp[2979]*kernel[1]+tmp[2980]*kernel[2]+tmp[3078]*kernel[3]+tmp[3079]*kernel[4]+tmp[3080]*kernel[5]+tmp[3178]*kernel[6]+tmp[3179]*kernel[7]+tmp[3180]*kernel[8];
				ans[3080]<=tmp[2979]*kernel[0]+tmp[2980]*kernel[1]+tmp[2981]*kernel[2]+tmp[3079]*kernel[3]+tmp[3080]*kernel[4]+tmp[3081]*kernel[5]+tmp[3179]*kernel[6]+tmp[3180]*kernel[7]+tmp[3181]*kernel[8];
				ans[3081]<=tmp[2980]*kernel[0]+tmp[2981]*kernel[1]+tmp[2982]*kernel[2]+tmp[3080]*kernel[3]+tmp[3081]*kernel[4]+tmp[3082]*kernel[5]+tmp[3180]*kernel[6]+tmp[3181]*kernel[7]+tmp[3182]*kernel[8];
				ans[3082]<=tmp[2981]*kernel[0]+tmp[2982]*kernel[1]+tmp[2983]*kernel[2]+tmp[3081]*kernel[3]+tmp[3082]*kernel[4]+tmp[3083]*kernel[5]+tmp[3181]*kernel[6]+tmp[3182]*kernel[7]+tmp[3183]*kernel[8];
				ans[3083]<=tmp[2982]*kernel[0]+tmp[2983]*kernel[1]+tmp[2984]*kernel[2]+tmp[3082]*kernel[3]+tmp[3083]*kernel[4]+tmp[3084]*kernel[5]+tmp[3182]*kernel[6]+tmp[3183]*kernel[7]+tmp[3184]*kernel[8];
				ans[3084]<=tmp[2983]*kernel[0]+tmp[2984]*kernel[1]+tmp[2985]*kernel[2]+tmp[3083]*kernel[3]+tmp[3084]*kernel[4]+tmp[3085]*kernel[5]+tmp[3183]*kernel[6]+tmp[3184]*kernel[7]+tmp[3185]*kernel[8];
				ans[3085]<=tmp[2984]*kernel[0]+tmp[2985]*kernel[1]+tmp[2986]*kernel[2]+tmp[3084]*kernel[3]+tmp[3085]*kernel[4]+tmp[3086]*kernel[5]+tmp[3184]*kernel[6]+tmp[3185]*kernel[7]+tmp[3186]*kernel[8];
				ans[3086]<=tmp[2985]*kernel[0]+tmp[2986]*kernel[1]+tmp[2987]*kernel[2]+tmp[3085]*kernel[3]+tmp[3086]*kernel[4]+tmp[3087]*kernel[5]+tmp[3185]*kernel[6]+tmp[3186]*kernel[7]+tmp[3187]*kernel[8];
				ans[3087]<=tmp[2986]*kernel[0]+tmp[2987]*kernel[1]+tmp[2988]*kernel[2]+tmp[3086]*kernel[3]+tmp[3087]*kernel[4]+tmp[3088]*kernel[5]+tmp[3186]*kernel[6]+tmp[3187]*kernel[7]+tmp[3188]*kernel[8];
				ans[3088]<=tmp[2987]*kernel[0]+tmp[2988]*kernel[1]+tmp[2989]*kernel[2]+tmp[3087]*kernel[3]+tmp[3088]*kernel[4]+tmp[3089]*kernel[5]+tmp[3187]*kernel[6]+tmp[3188]*kernel[7]+tmp[3189]*kernel[8];
				ans[3089]<=tmp[2988]*kernel[0]+tmp[2989]*kernel[1]+tmp[2990]*kernel[2]+tmp[3088]*kernel[3]+tmp[3089]*kernel[4]+tmp[3090]*kernel[5]+tmp[3188]*kernel[6]+tmp[3189]*kernel[7]+tmp[3190]*kernel[8];
				ans[3090]<=tmp[2989]*kernel[0]+tmp[2990]*kernel[1]+tmp[2991]*kernel[2]+tmp[3089]*kernel[3]+tmp[3090]*kernel[4]+tmp[3091]*kernel[5]+tmp[3189]*kernel[6]+tmp[3190]*kernel[7]+tmp[3191]*kernel[8];
				ans[3091]<=tmp[2990]*kernel[0]+tmp[2991]*kernel[1]+tmp[2992]*kernel[2]+tmp[3090]*kernel[3]+tmp[3091]*kernel[4]+tmp[3092]*kernel[5]+tmp[3190]*kernel[6]+tmp[3191]*kernel[7]+tmp[3192]*kernel[8];
				ans[3092]<=tmp[2991]*kernel[0]+tmp[2992]*kernel[1]+tmp[2993]*kernel[2]+tmp[3091]*kernel[3]+tmp[3092]*kernel[4]+tmp[3093]*kernel[5]+tmp[3191]*kernel[6]+tmp[3192]*kernel[7]+tmp[3193]*kernel[8];
				ans[3093]<=tmp[2992]*kernel[0]+tmp[2993]*kernel[1]+tmp[2994]*kernel[2]+tmp[3092]*kernel[3]+tmp[3093]*kernel[4]+tmp[3094]*kernel[5]+tmp[3192]*kernel[6]+tmp[3193]*kernel[7]+tmp[3194]*kernel[8];
				ans[3094]<=tmp[2993]*kernel[0]+tmp[2994]*kernel[1]+tmp[2995]*kernel[2]+tmp[3093]*kernel[3]+tmp[3094]*kernel[4]+tmp[3095]*kernel[5]+tmp[3193]*kernel[6]+tmp[3194]*kernel[7]+tmp[3195]*kernel[8];
				ans[3095]<=tmp[2994]*kernel[0]+tmp[2995]*kernel[1]+tmp[2996]*kernel[2]+tmp[3094]*kernel[3]+tmp[3095]*kernel[4]+tmp[3096]*kernel[5]+tmp[3194]*kernel[6]+tmp[3195]*kernel[7]+tmp[3196]*kernel[8];
				ans[3096]<=tmp[2995]*kernel[0]+tmp[2996]*kernel[1]+tmp[2997]*kernel[2]+tmp[3095]*kernel[3]+tmp[3096]*kernel[4]+tmp[3097]*kernel[5]+tmp[3195]*kernel[6]+tmp[3196]*kernel[7]+tmp[3197]*kernel[8];
				ans[3097]<=tmp[2996]*kernel[0]+tmp[2997]*kernel[1]+tmp[2998]*kernel[2]+tmp[3096]*kernel[3]+tmp[3097]*kernel[4]+tmp[3098]*kernel[5]+tmp[3196]*kernel[6]+tmp[3197]*kernel[7]+tmp[3198]*kernel[8];
				ans[3098]<=tmp[2997]*kernel[0]+tmp[2998]*kernel[1]+tmp[2999]*kernel[2]+tmp[3097]*kernel[3]+tmp[3098]*kernel[4]+tmp[3099]*kernel[5]+tmp[3197]*kernel[6]+tmp[3198]*kernel[7]+tmp[3199]*kernel[8];
				ans[3099]<=tmp[2998]*kernel[0]+tmp[2999]*kernel[1]+tmp[3098]*kernel[3]+tmp[3099]*kernel[4]+tmp[3198]*kernel[6]+tmp[3199]*kernel[7];
				ans[3100]<=tmp[3000]*kernel[1]+tmp[3001]*kernel[2]+tmp[3100]*kernel[4]+tmp[3101]*kernel[5]+tmp[3200]*kernel[7]+tmp[3201]*kernel[8];
				ans[3101]<=tmp[3000]*kernel[0]+tmp[3001]*kernel[1]+tmp[3002]*kernel[2]+tmp[3100]*kernel[3]+tmp[3101]*kernel[4]+tmp[3102]*kernel[5]+tmp[3200]*kernel[6]+tmp[3201]*kernel[7]+tmp[3202]*kernel[8];
				ans[3102]<=tmp[3001]*kernel[0]+tmp[3002]*kernel[1]+tmp[3003]*kernel[2]+tmp[3101]*kernel[3]+tmp[3102]*kernel[4]+tmp[3103]*kernel[5]+tmp[3201]*kernel[6]+tmp[3202]*kernel[7]+tmp[3203]*kernel[8];
				ans[3103]<=tmp[3002]*kernel[0]+tmp[3003]*kernel[1]+tmp[3004]*kernel[2]+tmp[3102]*kernel[3]+tmp[3103]*kernel[4]+tmp[3104]*kernel[5]+tmp[3202]*kernel[6]+tmp[3203]*kernel[7]+tmp[3204]*kernel[8];
				ans[3104]<=tmp[3003]*kernel[0]+tmp[3004]*kernel[1]+tmp[3005]*kernel[2]+tmp[3103]*kernel[3]+tmp[3104]*kernel[4]+tmp[3105]*kernel[5]+tmp[3203]*kernel[6]+tmp[3204]*kernel[7]+tmp[3205]*kernel[8];
				ans[3105]<=tmp[3004]*kernel[0]+tmp[3005]*kernel[1]+tmp[3006]*kernel[2]+tmp[3104]*kernel[3]+tmp[3105]*kernel[4]+tmp[3106]*kernel[5]+tmp[3204]*kernel[6]+tmp[3205]*kernel[7]+tmp[3206]*kernel[8];
				ans[3106]<=tmp[3005]*kernel[0]+tmp[3006]*kernel[1]+tmp[3007]*kernel[2]+tmp[3105]*kernel[3]+tmp[3106]*kernel[4]+tmp[3107]*kernel[5]+tmp[3205]*kernel[6]+tmp[3206]*kernel[7]+tmp[3207]*kernel[8];
				ans[3107]<=tmp[3006]*kernel[0]+tmp[3007]*kernel[1]+tmp[3008]*kernel[2]+tmp[3106]*kernel[3]+tmp[3107]*kernel[4]+tmp[3108]*kernel[5]+tmp[3206]*kernel[6]+tmp[3207]*kernel[7]+tmp[3208]*kernel[8];
				ans[3108]<=tmp[3007]*kernel[0]+tmp[3008]*kernel[1]+tmp[3009]*kernel[2]+tmp[3107]*kernel[3]+tmp[3108]*kernel[4]+tmp[3109]*kernel[5]+tmp[3207]*kernel[6]+tmp[3208]*kernel[7]+tmp[3209]*kernel[8];
				ans[3109]<=tmp[3008]*kernel[0]+tmp[3009]*kernel[1]+tmp[3010]*kernel[2]+tmp[3108]*kernel[3]+tmp[3109]*kernel[4]+tmp[3110]*kernel[5]+tmp[3208]*kernel[6]+tmp[3209]*kernel[7]+tmp[3210]*kernel[8];
				ans[3110]<=tmp[3009]*kernel[0]+tmp[3010]*kernel[1]+tmp[3011]*kernel[2]+tmp[3109]*kernel[3]+tmp[3110]*kernel[4]+tmp[3111]*kernel[5]+tmp[3209]*kernel[6]+tmp[3210]*kernel[7]+tmp[3211]*kernel[8];
				ans[3111]<=tmp[3010]*kernel[0]+tmp[3011]*kernel[1]+tmp[3012]*kernel[2]+tmp[3110]*kernel[3]+tmp[3111]*kernel[4]+tmp[3112]*kernel[5]+tmp[3210]*kernel[6]+tmp[3211]*kernel[7]+tmp[3212]*kernel[8];
				ans[3112]<=tmp[3011]*kernel[0]+tmp[3012]*kernel[1]+tmp[3013]*kernel[2]+tmp[3111]*kernel[3]+tmp[3112]*kernel[4]+tmp[3113]*kernel[5]+tmp[3211]*kernel[6]+tmp[3212]*kernel[7]+tmp[3213]*kernel[8];
				ans[3113]<=tmp[3012]*kernel[0]+tmp[3013]*kernel[1]+tmp[3014]*kernel[2]+tmp[3112]*kernel[3]+tmp[3113]*kernel[4]+tmp[3114]*kernel[5]+tmp[3212]*kernel[6]+tmp[3213]*kernel[7]+tmp[3214]*kernel[8];
				ans[3114]<=tmp[3013]*kernel[0]+tmp[3014]*kernel[1]+tmp[3015]*kernel[2]+tmp[3113]*kernel[3]+tmp[3114]*kernel[4]+tmp[3115]*kernel[5]+tmp[3213]*kernel[6]+tmp[3214]*kernel[7]+tmp[3215]*kernel[8];
				ans[3115]<=tmp[3014]*kernel[0]+tmp[3015]*kernel[1]+tmp[3016]*kernel[2]+tmp[3114]*kernel[3]+tmp[3115]*kernel[4]+tmp[3116]*kernel[5]+tmp[3214]*kernel[6]+tmp[3215]*kernel[7]+tmp[3216]*kernel[8];
				ans[3116]<=tmp[3015]*kernel[0]+tmp[3016]*kernel[1]+tmp[3017]*kernel[2]+tmp[3115]*kernel[3]+tmp[3116]*kernel[4]+tmp[3117]*kernel[5]+tmp[3215]*kernel[6]+tmp[3216]*kernel[7]+tmp[3217]*kernel[8];
				ans[3117]<=tmp[3016]*kernel[0]+tmp[3017]*kernel[1]+tmp[3018]*kernel[2]+tmp[3116]*kernel[3]+tmp[3117]*kernel[4]+tmp[3118]*kernel[5]+tmp[3216]*kernel[6]+tmp[3217]*kernel[7]+tmp[3218]*kernel[8];
				ans[3118]<=tmp[3017]*kernel[0]+tmp[3018]*kernel[1]+tmp[3019]*kernel[2]+tmp[3117]*kernel[3]+tmp[3118]*kernel[4]+tmp[3119]*kernel[5]+tmp[3217]*kernel[6]+tmp[3218]*kernel[7]+tmp[3219]*kernel[8];
				ans[3119]<=tmp[3018]*kernel[0]+tmp[3019]*kernel[1]+tmp[3020]*kernel[2]+tmp[3118]*kernel[3]+tmp[3119]*kernel[4]+tmp[3120]*kernel[5]+tmp[3218]*kernel[6]+tmp[3219]*kernel[7]+tmp[3220]*kernel[8];
				ans[3120]<=tmp[3019]*kernel[0]+tmp[3020]*kernel[1]+tmp[3021]*kernel[2]+tmp[3119]*kernel[3]+tmp[3120]*kernel[4]+tmp[3121]*kernel[5]+tmp[3219]*kernel[6]+tmp[3220]*kernel[7]+tmp[3221]*kernel[8];
				ans[3121]<=tmp[3020]*kernel[0]+tmp[3021]*kernel[1]+tmp[3022]*kernel[2]+tmp[3120]*kernel[3]+tmp[3121]*kernel[4]+tmp[3122]*kernel[5]+tmp[3220]*kernel[6]+tmp[3221]*kernel[7]+tmp[3222]*kernel[8];
				ans[3122]<=tmp[3021]*kernel[0]+tmp[3022]*kernel[1]+tmp[3023]*kernel[2]+tmp[3121]*kernel[3]+tmp[3122]*kernel[4]+tmp[3123]*kernel[5]+tmp[3221]*kernel[6]+tmp[3222]*kernel[7]+tmp[3223]*kernel[8];
				ans[3123]<=tmp[3022]*kernel[0]+tmp[3023]*kernel[1]+tmp[3024]*kernel[2]+tmp[3122]*kernel[3]+tmp[3123]*kernel[4]+tmp[3124]*kernel[5]+tmp[3222]*kernel[6]+tmp[3223]*kernel[7]+tmp[3224]*kernel[8];
				ans[3124]<=tmp[3023]*kernel[0]+tmp[3024]*kernel[1]+tmp[3025]*kernel[2]+tmp[3123]*kernel[3]+tmp[3124]*kernel[4]+tmp[3125]*kernel[5]+tmp[3223]*kernel[6]+tmp[3224]*kernel[7]+tmp[3225]*kernel[8];
				ans[3125]<=tmp[3024]*kernel[0]+tmp[3025]*kernel[1]+tmp[3026]*kernel[2]+tmp[3124]*kernel[3]+tmp[3125]*kernel[4]+tmp[3126]*kernel[5]+tmp[3224]*kernel[6]+tmp[3225]*kernel[7]+tmp[3226]*kernel[8];
				ans[3126]<=tmp[3025]*kernel[0]+tmp[3026]*kernel[1]+tmp[3027]*kernel[2]+tmp[3125]*kernel[3]+tmp[3126]*kernel[4]+tmp[3127]*kernel[5]+tmp[3225]*kernel[6]+tmp[3226]*kernel[7]+tmp[3227]*kernel[8];
				ans[3127]<=tmp[3026]*kernel[0]+tmp[3027]*kernel[1]+tmp[3028]*kernel[2]+tmp[3126]*kernel[3]+tmp[3127]*kernel[4]+tmp[3128]*kernel[5]+tmp[3226]*kernel[6]+tmp[3227]*kernel[7]+tmp[3228]*kernel[8];
				ans[3128]<=tmp[3027]*kernel[0]+tmp[3028]*kernel[1]+tmp[3029]*kernel[2]+tmp[3127]*kernel[3]+tmp[3128]*kernel[4]+tmp[3129]*kernel[5]+tmp[3227]*kernel[6]+tmp[3228]*kernel[7]+tmp[3229]*kernel[8];
				ans[3129]<=tmp[3028]*kernel[0]+tmp[3029]*kernel[1]+tmp[3030]*kernel[2]+tmp[3128]*kernel[3]+tmp[3129]*kernel[4]+tmp[3130]*kernel[5]+tmp[3228]*kernel[6]+tmp[3229]*kernel[7]+tmp[3230]*kernel[8];
				ans[3130]<=tmp[3029]*kernel[0]+tmp[3030]*kernel[1]+tmp[3031]*kernel[2]+tmp[3129]*kernel[3]+tmp[3130]*kernel[4]+tmp[3131]*kernel[5]+tmp[3229]*kernel[6]+tmp[3230]*kernel[7]+tmp[3231]*kernel[8];
				ans[3131]<=tmp[3030]*kernel[0]+tmp[3031]*kernel[1]+tmp[3032]*kernel[2]+tmp[3130]*kernel[3]+tmp[3131]*kernel[4]+tmp[3132]*kernel[5]+tmp[3230]*kernel[6]+tmp[3231]*kernel[7]+tmp[3232]*kernel[8];
				ans[3132]<=tmp[3031]*kernel[0]+tmp[3032]*kernel[1]+tmp[3033]*kernel[2]+tmp[3131]*kernel[3]+tmp[3132]*kernel[4]+tmp[3133]*kernel[5]+tmp[3231]*kernel[6]+tmp[3232]*kernel[7]+tmp[3233]*kernel[8];
				ans[3133]<=tmp[3032]*kernel[0]+tmp[3033]*kernel[1]+tmp[3034]*kernel[2]+tmp[3132]*kernel[3]+tmp[3133]*kernel[4]+tmp[3134]*kernel[5]+tmp[3232]*kernel[6]+tmp[3233]*kernel[7]+tmp[3234]*kernel[8];
				ans[3134]<=tmp[3033]*kernel[0]+tmp[3034]*kernel[1]+tmp[3035]*kernel[2]+tmp[3133]*kernel[3]+tmp[3134]*kernel[4]+tmp[3135]*kernel[5]+tmp[3233]*kernel[6]+tmp[3234]*kernel[7]+tmp[3235]*kernel[8];
				ans[3135]<=tmp[3034]*kernel[0]+tmp[3035]*kernel[1]+tmp[3036]*kernel[2]+tmp[3134]*kernel[3]+tmp[3135]*kernel[4]+tmp[3136]*kernel[5]+tmp[3234]*kernel[6]+tmp[3235]*kernel[7]+tmp[3236]*kernel[8];
				ans[3136]<=tmp[3035]*kernel[0]+tmp[3036]*kernel[1]+tmp[3037]*kernel[2]+tmp[3135]*kernel[3]+tmp[3136]*kernel[4]+tmp[3137]*kernel[5]+tmp[3235]*kernel[6]+tmp[3236]*kernel[7]+tmp[3237]*kernel[8];
				ans[3137]<=tmp[3036]*kernel[0]+tmp[3037]*kernel[1]+tmp[3038]*kernel[2]+tmp[3136]*kernel[3]+tmp[3137]*kernel[4]+tmp[3138]*kernel[5]+tmp[3236]*kernel[6]+tmp[3237]*kernel[7]+tmp[3238]*kernel[8];
				ans[3138]<=tmp[3037]*kernel[0]+tmp[3038]*kernel[1]+tmp[3039]*kernel[2]+tmp[3137]*kernel[3]+tmp[3138]*kernel[4]+tmp[3139]*kernel[5]+tmp[3237]*kernel[6]+tmp[3238]*kernel[7]+tmp[3239]*kernel[8];
				ans[3139]<=tmp[3038]*kernel[0]+tmp[3039]*kernel[1]+tmp[3040]*kernel[2]+tmp[3138]*kernel[3]+tmp[3139]*kernel[4]+tmp[3140]*kernel[5]+tmp[3238]*kernel[6]+tmp[3239]*kernel[7]+tmp[3240]*kernel[8];
				ans[3140]<=tmp[3039]*kernel[0]+tmp[3040]*kernel[1]+tmp[3041]*kernel[2]+tmp[3139]*kernel[3]+tmp[3140]*kernel[4]+tmp[3141]*kernel[5]+tmp[3239]*kernel[6]+tmp[3240]*kernel[7]+tmp[3241]*kernel[8];
				ans[3141]<=tmp[3040]*kernel[0]+tmp[3041]*kernel[1]+tmp[3042]*kernel[2]+tmp[3140]*kernel[3]+tmp[3141]*kernel[4]+tmp[3142]*kernel[5]+tmp[3240]*kernel[6]+tmp[3241]*kernel[7]+tmp[3242]*kernel[8];
				ans[3142]<=tmp[3041]*kernel[0]+tmp[3042]*kernel[1]+tmp[3043]*kernel[2]+tmp[3141]*kernel[3]+tmp[3142]*kernel[4]+tmp[3143]*kernel[5]+tmp[3241]*kernel[6]+tmp[3242]*kernel[7]+tmp[3243]*kernel[8];
				ans[3143]<=tmp[3042]*kernel[0]+tmp[3043]*kernel[1]+tmp[3044]*kernel[2]+tmp[3142]*kernel[3]+tmp[3143]*kernel[4]+tmp[3144]*kernel[5]+tmp[3242]*kernel[6]+tmp[3243]*kernel[7]+tmp[3244]*kernel[8];
				ans[3144]<=tmp[3043]*kernel[0]+tmp[3044]*kernel[1]+tmp[3045]*kernel[2]+tmp[3143]*kernel[3]+tmp[3144]*kernel[4]+tmp[3145]*kernel[5]+tmp[3243]*kernel[6]+tmp[3244]*kernel[7]+tmp[3245]*kernel[8];
				ans[3145]<=tmp[3044]*kernel[0]+tmp[3045]*kernel[1]+tmp[3046]*kernel[2]+tmp[3144]*kernel[3]+tmp[3145]*kernel[4]+tmp[3146]*kernel[5]+tmp[3244]*kernel[6]+tmp[3245]*kernel[7]+tmp[3246]*kernel[8];
				ans[3146]<=tmp[3045]*kernel[0]+tmp[3046]*kernel[1]+tmp[3047]*kernel[2]+tmp[3145]*kernel[3]+tmp[3146]*kernel[4]+tmp[3147]*kernel[5]+tmp[3245]*kernel[6]+tmp[3246]*kernel[7]+tmp[3247]*kernel[8];
				ans[3147]<=tmp[3046]*kernel[0]+tmp[3047]*kernel[1]+tmp[3048]*kernel[2]+tmp[3146]*kernel[3]+tmp[3147]*kernel[4]+tmp[3148]*kernel[5]+tmp[3246]*kernel[6]+tmp[3247]*kernel[7]+tmp[3248]*kernel[8];
				ans[3148]<=tmp[3047]*kernel[0]+tmp[3048]*kernel[1]+tmp[3049]*kernel[2]+tmp[3147]*kernel[3]+tmp[3148]*kernel[4]+tmp[3149]*kernel[5]+tmp[3247]*kernel[6]+tmp[3248]*kernel[7]+tmp[3249]*kernel[8];
				ans[3149]<=tmp[3048]*kernel[0]+tmp[3049]*kernel[1]+tmp[3050]*kernel[2]+tmp[3148]*kernel[3]+tmp[3149]*kernel[4]+tmp[3150]*kernel[5]+tmp[3248]*kernel[6]+tmp[3249]*kernel[7]+tmp[3250]*kernel[8];
				ans[3150]<=tmp[3049]*kernel[0]+tmp[3050]*kernel[1]+tmp[3051]*kernel[2]+tmp[3149]*kernel[3]+tmp[3150]*kernel[4]+tmp[3151]*kernel[5]+tmp[3249]*kernel[6]+tmp[3250]*kernel[7]+tmp[3251]*kernel[8];
				ans[3151]<=tmp[3050]*kernel[0]+tmp[3051]*kernel[1]+tmp[3052]*kernel[2]+tmp[3150]*kernel[3]+tmp[3151]*kernel[4]+tmp[3152]*kernel[5]+tmp[3250]*kernel[6]+tmp[3251]*kernel[7]+tmp[3252]*kernel[8];
				ans[3152]<=tmp[3051]*kernel[0]+tmp[3052]*kernel[1]+tmp[3053]*kernel[2]+tmp[3151]*kernel[3]+tmp[3152]*kernel[4]+tmp[3153]*kernel[5]+tmp[3251]*kernel[6]+tmp[3252]*kernel[7]+tmp[3253]*kernel[8];
				ans[3153]<=tmp[3052]*kernel[0]+tmp[3053]*kernel[1]+tmp[3054]*kernel[2]+tmp[3152]*kernel[3]+tmp[3153]*kernel[4]+tmp[3154]*kernel[5]+tmp[3252]*kernel[6]+tmp[3253]*kernel[7]+tmp[3254]*kernel[8];
				ans[3154]<=tmp[3053]*kernel[0]+tmp[3054]*kernel[1]+tmp[3055]*kernel[2]+tmp[3153]*kernel[3]+tmp[3154]*kernel[4]+tmp[3155]*kernel[5]+tmp[3253]*kernel[6]+tmp[3254]*kernel[7]+tmp[3255]*kernel[8];
				ans[3155]<=tmp[3054]*kernel[0]+tmp[3055]*kernel[1]+tmp[3056]*kernel[2]+tmp[3154]*kernel[3]+tmp[3155]*kernel[4]+tmp[3156]*kernel[5]+tmp[3254]*kernel[6]+tmp[3255]*kernel[7]+tmp[3256]*kernel[8];
				ans[3156]<=tmp[3055]*kernel[0]+tmp[3056]*kernel[1]+tmp[3057]*kernel[2]+tmp[3155]*kernel[3]+tmp[3156]*kernel[4]+tmp[3157]*kernel[5]+tmp[3255]*kernel[6]+tmp[3256]*kernel[7]+tmp[3257]*kernel[8];
				ans[3157]<=tmp[3056]*kernel[0]+tmp[3057]*kernel[1]+tmp[3058]*kernel[2]+tmp[3156]*kernel[3]+tmp[3157]*kernel[4]+tmp[3158]*kernel[5]+tmp[3256]*kernel[6]+tmp[3257]*kernel[7]+tmp[3258]*kernel[8];
				ans[3158]<=tmp[3057]*kernel[0]+tmp[3058]*kernel[1]+tmp[3059]*kernel[2]+tmp[3157]*kernel[3]+tmp[3158]*kernel[4]+tmp[3159]*kernel[5]+tmp[3257]*kernel[6]+tmp[3258]*kernel[7]+tmp[3259]*kernel[8];
				ans[3159]<=tmp[3058]*kernel[0]+tmp[3059]*kernel[1]+tmp[3060]*kernel[2]+tmp[3158]*kernel[3]+tmp[3159]*kernel[4]+tmp[3160]*kernel[5]+tmp[3258]*kernel[6]+tmp[3259]*kernel[7]+tmp[3260]*kernel[8];
				ans[3160]<=tmp[3059]*kernel[0]+tmp[3060]*kernel[1]+tmp[3061]*kernel[2]+tmp[3159]*kernel[3]+tmp[3160]*kernel[4]+tmp[3161]*kernel[5]+tmp[3259]*kernel[6]+tmp[3260]*kernel[7]+tmp[3261]*kernel[8];
				ans[3161]<=tmp[3060]*kernel[0]+tmp[3061]*kernel[1]+tmp[3062]*kernel[2]+tmp[3160]*kernel[3]+tmp[3161]*kernel[4]+tmp[3162]*kernel[5]+tmp[3260]*kernel[6]+tmp[3261]*kernel[7]+tmp[3262]*kernel[8];
				ans[3162]<=tmp[3061]*kernel[0]+tmp[3062]*kernel[1]+tmp[3063]*kernel[2]+tmp[3161]*kernel[3]+tmp[3162]*kernel[4]+tmp[3163]*kernel[5]+tmp[3261]*kernel[6]+tmp[3262]*kernel[7]+tmp[3263]*kernel[8];
				ans[3163]<=tmp[3062]*kernel[0]+tmp[3063]*kernel[1]+tmp[3064]*kernel[2]+tmp[3162]*kernel[3]+tmp[3163]*kernel[4]+tmp[3164]*kernel[5]+tmp[3262]*kernel[6]+tmp[3263]*kernel[7]+tmp[3264]*kernel[8];
				ans[3164]<=tmp[3063]*kernel[0]+tmp[3064]*kernel[1]+tmp[3065]*kernel[2]+tmp[3163]*kernel[3]+tmp[3164]*kernel[4]+tmp[3165]*kernel[5]+tmp[3263]*kernel[6]+tmp[3264]*kernel[7]+tmp[3265]*kernel[8];
				ans[3165]<=tmp[3064]*kernel[0]+tmp[3065]*kernel[1]+tmp[3066]*kernel[2]+tmp[3164]*kernel[3]+tmp[3165]*kernel[4]+tmp[3166]*kernel[5]+tmp[3264]*kernel[6]+tmp[3265]*kernel[7]+tmp[3266]*kernel[8];
				ans[3166]<=tmp[3065]*kernel[0]+tmp[3066]*kernel[1]+tmp[3067]*kernel[2]+tmp[3165]*kernel[3]+tmp[3166]*kernel[4]+tmp[3167]*kernel[5]+tmp[3265]*kernel[6]+tmp[3266]*kernel[7]+tmp[3267]*kernel[8];
				ans[3167]<=tmp[3066]*kernel[0]+tmp[3067]*kernel[1]+tmp[3068]*kernel[2]+tmp[3166]*kernel[3]+tmp[3167]*kernel[4]+tmp[3168]*kernel[5]+tmp[3266]*kernel[6]+tmp[3267]*kernel[7]+tmp[3268]*kernel[8];
				ans[3168]<=tmp[3067]*kernel[0]+tmp[3068]*kernel[1]+tmp[3069]*kernel[2]+tmp[3167]*kernel[3]+tmp[3168]*kernel[4]+tmp[3169]*kernel[5]+tmp[3267]*kernel[6]+tmp[3268]*kernel[7]+tmp[3269]*kernel[8];
				ans[3169]<=tmp[3068]*kernel[0]+tmp[3069]*kernel[1]+tmp[3070]*kernel[2]+tmp[3168]*kernel[3]+tmp[3169]*kernel[4]+tmp[3170]*kernel[5]+tmp[3268]*kernel[6]+tmp[3269]*kernel[7]+tmp[3270]*kernel[8];
				ans[3170]<=tmp[3069]*kernel[0]+tmp[3070]*kernel[1]+tmp[3071]*kernel[2]+tmp[3169]*kernel[3]+tmp[3170]*kernel[4]+tmp[3171]*kernel[5]+tmp[3269]*kernel[6]+tmp[3270]*kernel[7]+tmp[3271]*kernel[8];
				ans[3171]<=tmp[3070]*kernel[0]+tmp[3071]*kernel[1]+tmp[3072]*kernel[2]+tmp[3170]*kernel[3]+tmp[3171]*kernel[4]+tmp[3172]*kernel[5]+tmp[3270]*kernel[6]+tmp[3271]*kernel[7]+tmp[3272]*kernel[8];
				ans[3172]<=tmp[3071]*kernel[0]+tmp[3072]*kernel[1]+tmp[3073]*kernel[2]+tmp[3171]*kernel[3]+tmp[3172]*kernel[4]+tmp[3173]*kernel[5]+tmp[3271]*kernel[6]+tmp[3272]*kernel[7]+tmp[3273]*kernel[8];
				ans[3173]<=tmp[3072]*kernel[0]+tmp[3073]*kernel[1]+tmp[3074]*kernel[2]+tmp[3172]*kernel[3]+tmp[3173]*kernel[4]+tmp[3174]*kernel[5]+tmp[3272]*kernel[6]+tmp[3273]*kernel[7]+tmp[3274]*kernel[8];
				ans[3174]<=tmp[3073]*kernel[0]+tmp[3074]*kernel[1]+tmp[3075]*kernel[2]+tmp[3173]*kernel[3]+tmp[3174]*kernel[4]+tmp[3175]*kernel[5]+tmp[3273]*kernel[6]+tmp[3274]*kernel[7]+tmp[3275]*kernel[8];
				ans[3175]<=tmp[3074]*kernel[0]+tmp[3075]*kernel[1]+tmp[3076]*kernel[2]+tmp[3174]*kernel[3]+tmp[3175]*kernel[4]+tmp[3176]*kernel[5]+tmp[3274]*kernel[6]+tmp[3275]*kernel[7]+tmp[3276]*kernel[8];
				ans[3176]<=tmp[3075]*kernel[0]+tmp[3076]*kernel[1]+tmp[3077]*kernel[2]+tmp[3175]*kernel[3]+tmp[3176]*kernel[4]+tmp[3177]*kernel[5]+tmp[3275]*kernel[6]+tmp[3276]*kernel[7]+tmp[3277]*kernel[8];
				ans[3177]<=tmp[3076]*kernel[0]+tmp[3077]*kernel[1]+tmp[3078]*kernel[2]+tmp[3176]*kernel[3]+tmp[3177]*kernel[4]+tmp[3178]*kernel[5]+tmp[3276]*kernel[6]+tmp[3277]*kernel[7]+tmp[3278]*kernel[8];
				ans[3178]<=tmp[3077]*kernel[0]+tmp[3078]*kernel[1]+tmp[3079]*kernel[2]+tmp[3177]*kernel[3]+tmp[3178]*kernel[4]+tmp[3179]*kernel[5]+tmp[3277]*kernel[6]+tmp[3278]*kernel[7]+tmp[3279]*kernel[8];
				ans[3179]<=tmp[3078]*kernel[0]+tmp[3079]*kernel[1]+tmp[3080]*kernel[2]+tmp[3178]*kernel[3]+tmp[3179]*kernel[4]+tmp[3180]*kernel[5]+tmp[3278]*kernel[6]+tmp[3279]*kernel[7]+tmp[3280]*kernel[8];
				ans[3180]<=tmp[3079]*kernel[0]+tmp[3080]*kernel[1]+tmp[3081]*kernel[2]+tmp[3179]*kernel[3]+tmp[3180]*kernel[4]+tmp[3181]*kernel[5]+tmp[3279]*kernel[6]+tmp[3280]*kernel[7]+tmp[3281]*kernel[8];
				ans[3181]<=tmp[3080]*kernel[0]+tmp[3081]*kernel[1]+tmp[3082]*kernel[2]+tmp[3180]*kernel[3]+tmp[3181]*kernel[4]+tmp[3182]*kernel[5]+tmp[3280]*kernel[6]+tmp[3281]*kernel[7]+tmp[3282]*kernel[8];
				ans[3182]<=tmp[3081]*kernel[0]+tmp[3082]*kernel[1]+tmp[3083]*kernel[2]+tmp[3181]*kernel[3]+tmp[3182]*kernel[4]+tmp[3183]*kernel[5]+tmp[3281]*kernel[6]+tmp[3282]*kernel[7]+tmp[3283]*kernel[8];
				ans[3183]<=tmp[3082]*kernel[0]+tmp[3083]*kernel[1]+tmp[3084]*kernel[2]+tmp[3182]*kernel[3]+tmp[3183]*kernel[4]+tmp[3184]*kernel[5]+tmp[3282]*kernel[6]+tmp[3283]*kernel[7]+tmp[3284]*kernel[8];
				ans[3184]<=tmp[3083]*kernel[0]+tmp[3084]*kernel[1]+tmp[3085]*kernel[2]+tmp[3183]*kernel[3]+tmp[3184]*kernel[4]+tmp[3185]*kernel[5]+tmp[3283]*kernel[6]+tmp[3284]*kernel[7]+tmp[3285]*kernel[8];
				ans[3185]<=tmp[3084]*kernel[0]+tmp[3085]*kernel[1]+tmp[3086]*kernel[2]+tmp[3184]*kernel[3]+tmp[3185]*kernel[4]+tmp[3186]*kernel[5]+tmp[3284]*kernel[6]+tmp[3285]*kernel[7]+tmp[3286]*kernel[8];
				ans[3186]<=tmp[3085]*kernel[0]+tmp[3086]*kernel[1]+tmp[3087]*kernel[2]+tmp[3185]*kernel[3]+tmp[3186]*kernel[4]+tmp[3187]*kernel[5]+tmp[3285]*kernel[6]+tmp[3286]*kernel[7]+tmp[3287]*kernel[8];
				ans[3187]<=tmp[3086]*kernel[0]+tmp[3087]*kernel[1]+tmp[3088]*kernel[2]+tmp[3186]*kernel[3]+tmp[3187]*kernel[4]+tmp[3188]*kernel[5]+tmp[3286]*kernel[6]+tmp[3287]*kernel[7]+tmp[3288]*kernel[8];
				ans[3188]<=tmp[3087]*kernel[0]+tmp[3088]*kernel[1]+tmp[3089]*kernel[2]+tmp[3187]*kernel[3]+tmp[3188]*kernel[4]+tmp[3189]*kernel[5]+tmp[3287]*kernel[6]+tmp[3288]*kernel[7]+tmp[3289]*kernel[8];
				ans[3189]<=tmp[3088]*kernel[0]+tmp[3089]*kernel[1]+tmp[3090]*kernel[2]+tmp[3188]*kernel[3]+tmp[3189]*kernel[4]+tmp[3190]*kernel[5]+tmp[3288]*kernel[6]+tmp[3289]*kernel[7]+tmp[3290]*kernel[8];
				ans[3190]<=tmp[3089]*kernel[0]+tmp[3090]*kernel[1]+tmp[3091]*kernel[2]+tmp[3189]*kernel[3]+tmp[3190]*kernel[4]+tmp[3191]*kernel[5]+tmp[3289]*kernel[6]+tmp[3290]*kernel[7]+tmp[3291]*kernel[8];
				ans[3191]<=tmp[3090]*kernel[0]+tmp[3091]*kernel[1]+tmp[3092]*kernel[2]+tmp[3190]*kernel[3]+tmp[3191]*kernel[4]+tmp[3192]*kernel[5]+tmp[3290]*kernel[6]+tmp[3291]*kernel[7]+tmp[3292]*kernel[8];
				ans[3192]<=tmp[3091]*kernel[0]+tmp[3092]*kernel[1]+tmp[3093]*kernel[2]+tmp[3191]*kernel[3]+tmp[3192]*kernel[4]+tmp[3193]*kernel[5]+tmp[3291]*kernel[6]+tmp[3292]*kernel[7]+tmp[3293]*kernel[8];
				ans[3193]<=tmp[3092]*kernel[0]+tmp[3093]*kernel[1]+tmp[3094]*kernel[2]+tmp[3192]*kernel[3]+tmp[3193]*kernel[4]+tmp[3194]*kernel[5]+tmp[3292]*kernel[6]+tmp[3293]*kernel[7]+tmp[3294]*kernel[8];
				ans[3194]<=tmp[3093]*kernel[0]+tmp[3094]*kernel[1]+tmp[3095]*kernel[2]+tmp[3193]*kernel[3]+tmp[3194]*kernel[4]+tmp[3195]*kernel[5]+tmp[3293]*kernel[6]+tmp[3294]*kernel[7]+tmp[3295]*kernel[8];
				ans[3195]<=tmp[3094]*kernel[0]+tmp[3095]*kernel[1]+tmp[3096]*kernel[2]+tmp[3194]*kernel[3]+tmp[3195]*kernel[4]+tmp[3196]*kernel[5]+tmp[3294]*kernel[6]+tmp[3295]*kernel[7]+tmp[3296]*kernel[8];
				ans[3196]<=tmp[3095]*kernel[0]+tmp[3096]*kernel[1]+tmp[3097]*kernel[2]+tmp[3195]*kernel[3]+tmp[3196]*kernel[4]+tmp[3197]*kernel[5]+tmp[3295]*kernel[6]+tmp[3296]*kernel[7]+tmp[3297]*kernel[8];
				ans[3197]<=tmp[3096]*kernel[0]+tmp[3097]*kernel[1]+tmp[3098]*kernel[2]+tmp[3196]*kernel[3]+tmp[3197]*kernel[4]+tmp[3198]*kernel[5]+tmp[3296]*kernel[6]+tmp[3297]*kernel[7]+tmp[3298]*kernel[8];
				ans[3198]<=tmp[3097]*kernel[0]+tmp[3098]*kernel[1]+tmp[3099]*kernel[2]+tmp[3197]*kernel[3]+tmp[3198]*kernel[4]+tmp[3199]*kernel[5]+tmp[3297]*kernel[6]+tmp[3298]*kernel[7]+tmp[3299]*kernel[8];
				ans[3199]<=tmp[3098]*kernel[0]+tmp[3099]*kernel[1]+tmp[3198]*kernel[3]+tmp[3199]*kernel[4]+tmp[3298]*kernel[6]+tmp[3299]*kernel[7];
				ans[3200]<=tmp[3100]*kernel[1]+tmp[3101]*kernel[2]+tmp[3200]*kernel[4]+tmp[3201]*kernel[5]+tmp[3300]*kernel[7]+tmp[3301]*kernel[8];
				ans[3201]<=tmp[3100]*kernel[0]+tmp[3101]*kernel[1]+tmp[3102]*kernel[2]+tmp[3200]*kernel[3]+tmp[3201]*kernel[4]+tmp[3202]*kernel[5]+tmp[3300]*kernel[6]+tmp[3301]*kernel[7]+tmp[3302]*kernel[8];
				ans[3202]<=tmp[3101]*kernel[0]+tmp[3102]*kernel[1]+tmp[3103]*kernel[2]+tmp[3201]*kernel[3]+tmp[3202]*kernel[4]+tmp[3203]*kernel[5]+tmp[3301]*kernel[6]+tmp[3302]*kernel[7]+tmp[3303]*kernel[8];
				ans[3203]<=tmp[3102]*kernel[0]+tmp[3103]*kernel[1]+tmp[3104]*kernel[2]+tmp[3202]*kernel[3]+tmp[3203]*kernel[4]+tmp[3204]*kernel[5]+tmp[3302]*kernel[6]+tmp[3303]*kernel[7]+tmp[3304]*kernel[8];
				ans[3204]<=tmp[3103]*kernel[0]+tmp[3104]*kernel[1]+tmp[3105]*kernel[2]+tmp[3203]*kernel[3]+tmp[3204]*kernel[4]+tmp[3205]*kernel[5]+tmp[3303]*kernel[6]+tmp[3304]*kernel[7]+tmp[3305]*kernel[8];
				ans[3205]<=tmp[3104]*kernel[0]+tmp[3105]*kernel[1]+tmp[3106]*kernel[2]+tmp[3204]*kernel[3]+tmp[3205]*kernel[4]+tmp[3206]*kernel[5]+tmp[3304]*kernel[6]+tmp[3305]*kernel[7]+tmp[3306]*kernel[8];
				ans[3206]<=tmp[3105]*kernel[0]+tmp[3106]*kernel[1]+tmp[3107]*kernel[2]+tmp[3205]*kernel[3]+tmp[3206]*kernel[4]+tmp[3207]*kernel[5]+tmp[3305]*kernel[6]+tmp[3306]*kernel[7]+tmp[3307]*kernel[8];
				ans[3207]<=tmp[3106]*kernel[0]+tmp[3107]*kernel[1]+tmp[3108]*kernel[2]+tmp[3206]*kernel[3]+tmp[3207]*kernel[4]+tmp[3208]*kernel[5]+tmp[3306]*kernel[6]+tmp[3307]*kernel[7]+tmp[3308]*kernel[8];
				ans[3208]<=tmp[3107]*kernel[0]+tmp[3108]*kernel[1]+tmp[3109]*kernel[2]+tmp[3207]*kernel[3]+tmp[3208]*kernel[4]+tmp[3209]*kernel[5]+tmp[3307]*kernel[6]+tmp[3308]*kernel[7]+tmp[3309]*kernel[8];
				ans[3209]<=tmp[3108]*kernel[0]+tmp[3109]*kernel[1]+tmp[3110]*kernel[2]+tmp[3208]*kernel[3]+tmp[3209]*kernel[4]+tmp[3210]*kernel[5]+tmp[3308]*kernel[6]+tmp[3309]*kernel[7]+tmp[3310]*kernel[8];
				ans[3210]<=tmp[3109]*kernel[0]+tmp[3110]*kernel[1]+tmp[3111]*kernel[2]+tmp[3209]*kernel[3]+tmp[3210]*kernel[4]+tmp[3211]*kernel[5]+tmp[3309]*kernel[6]+tmp[3310]*kernel[7]+tmp[3311]*kernel[8];
				ans[3211]<=tmp[3110]*kernel[0]+tmp[3111]*kernel[1]+tmp[3112]*kernel[2]+tmp[3210]*kernel[3]+tmp[3211]*kernel[4]+tmp[3212]*kernel[5]+tmp[3310]*kernel[6]+tmp[3311]*kernel[7]+tmp[3312]*kernel[8];
				ans[3212]<=tmp[3111]*kernel[0]+tmp[3112]*kernel[1]+tmp[3113]*kernel[2]+tmp[3211]*kernel[3]+tmp[3212]*kernel[4]+tmp[3213]*kernel[5]+tmp[3311]*kernel[6]+tmp[3312]*kernel[7]+tmp[3313]*kernel[8];
				ans[3213]<=tmp[3112]*kernel[0]+tmp[3113]*kernel[1]+tmp[3114]*kernel[2]+tmp[3212]*kernel[3]+tmp[3213]*kernel[4]+tmp[3214]*kernel[5]+tmp[3312]*kernel[6]+tmp[3313]*kernel[7]+tmp[3314]*kernel[8];
				ans[3214]<=tmp[3113]*kernel[0]+tmp[3114]*kernel[1]+tmp[3115]*kernel[2]+tmp[3213]*kernel[3]+tmp[3214]*kernel[4]+tmp[3215]*kernel[5]+tmp[3313]*kernel[6]+tmp[3314]*kernel[7]+tmp[3315]*kernel[8];
				ans[3215]<=tmp[3114]*kernel[0]+tmp[3115]*kernel[1]+tmp[3116]*kernel[2]+tmp[3214]*kernel[3]+tmp[3215]*kernel[4]+tmp[3216]*kernel[5]+tmp[3314]*kernel[6]+tmp[3315]*kernel[7]+tmp[3316]*kernel[8];
				ans[3216]<=tmp[3115]*kernel[0]+tmp[3116]*kernel[1]+tmp[3117]*kernel[2]+tmp[3215]*kernel[3]+tmp[3216]*kernel[4]+tmp[3217]*kernel[5]+tmp[3315]*kernel[6]+tmp[3316]*kernel[7]+tmp[3317]*kernel[8];
				ans[3217]<=tmp[3116]*kernel[0]+tmp[3117]*kernel[1]+tmp[3118]*kernel[2]+tmp[3216]*kernel[3]+tmp[3217]*kernel[4]+tmp[3218]*kernel[5]+tmp[3316]*kernel[6]+tmp[3317]*kernel[7]+tmp[3318]*kernel[8];
				ans[3218]<=tmp[3117]*kernel[0]+tmp[3118]*kernel[1]+tmp[3119]*kernel[2]+tmp[3217]*kernel[3]+tmp[3218]*kernel[4]+tmp[3219]*kernel[5]+tmp[3317]*kernel[6]+tmp[3318]*kernel[7]+tmp[3319]*kernel[8];
				ans[3219]<=tmp[3118]*kernel[0]+tmp[3119]*kernel[1]+tmp[3120]*kernel[2]+tmp[3218]*kernel[3]+tmp[3219]*kernel[4]+tmp[3220]*kernel[5]+tmp[3318]*kernel[6]+tmp[3319]*kernel[7]+tmp[3320]*kernel[8];
				ans[3220]<=tmp[3119]*kernel[0]+tmp[3120]*kernel[1]+tmp[3121]*kernel[2]+tmp[3219]*kernel[3]+tmp[3220]*kernel[4]+tmp[3221]*kernel[5]+tmp[3319]*kernel[6]+tmp[3320]*kernel[7]+tmp[3321]*kernel[8];
				ans[3221]<=tmp[3120]*kernel[0]+tmp[3121]*kernel[1]+tmp[3122]*kernel[2]+tmp[3220]*kernel[3]+tmp[3221]*kernel[4]+tmp[3222]*kernel[5]+tmp[3320]*kernel[6]+tmp[3321]*kernel[7]+tmp[3322]*kernel[8];
				ans[3222]<=tmp[3121]*kernel[0]+tmp[3122]*kernel[1]+tmp[3123]*kernel[2]+tmp[3221]*kernel[3]+tmp[3222]*kernel[4]+tmp[3223]*kernel[5]+tmp[3321]*kernel[6]+tmp[3322]*kernel[7]+tmp[3323]*kernel[8];
				ans[3223]<=tmp[3122]*kernel[0]+tmp[3123]*kernel[1]+tmp[3124]*kernel[2]+tmp[3222]*kernel[3]+tmp[3223]*kernel[4]+tmp[3224]*kernel[5]+tmp[3322]*kernel[6]+tmp[3323]*kernel[7]+tmp[3324]*kernel[8];
				ans[3224]<=tmp[3123]*kernel[0]+tmp[3124]*kernel[1]+tmp[3125]*kernel[2]+tmp[3223]*kernel[3]+tmp[3224]*kernel[4]+tmp[3225]*kernel[5]+tmp[3323]*kernel[6]+tmp[3324]*kernel[7]+tmp[3325]*kernel[8];
				ans[3225]<=tmp[3124]*kernel[0]+tmp[3125]*kernel[1]+tmp[3126]*kernel[2]+tmp[3224]*kernel[3]+tmp[3225]*kernel[4]+tmp[3226]*kernel[5]+tmp[3324]*kernel[6]+tmp[3325]*kernel[7]+tmp[3326]*kernel[8];
				ans[3226]<=tmp[3125]*kernel[0]+tmp[3126]*kernel[1]+tmp[3127]*kernel[2]+tmp[3225]*kernel[3]+tmp[3226]*kernel[4]+tmp[3227]*kernel[5]+tmp[3325]*kernel[6]+tmp[3326]*kernel[7]+tmp[3327]*kernel[8];
				ans[3227]<=tmp[3126]*kernel[0]+tmp[3127]*kernel[1]+tmp[3128]*kernel[2]+tmp[3226]*kernel[3]+tmp[3227]*kernel[4]+tmp[3228]*kernel[5]+tmp[3326]*kernel[6]+tmp[3327]*kernel[7]+tmp[3328]*kernel[8];
				ans[3228]<=tmp[3127]*kernel[0]+tmp[3128]*kernel[1]+tmp[3129]*kernel[2]+tmp[3227]*kernel[3]+tmp[3228]*kernel[4]+tmp[3229]*kernel[5]+tmp[3327]*kernel[6]+tmp[3328]*kernel[7]+tmp[3329]*kernel[8];
				ans[3229]<=tmp[3128]*kernel[0]+tmp[3129]*kernel[1]+tmp[3130]*kernel[2]+tmp[3228]*kernel[3]+tmp[3229]*kernel[4]+tmp[3230]*kernel[5]+tmp[3328]*kernel[6]+tmp[3329]*kernel[7]+tmp[3330]*kernel[8];
				ans[3230]<=tmp[3129]*kernel[0]+tmp[3130]*kernel[1]+tmp[3131]*kernel[2]+tmp[3229]*kernel[3]+tmp[3230]*kernel[4]+tmp[3231]*kernel[5]+tmp[3329]*kernel[6]+tmp[3330]*kernel[7]+tmp[3331]*kernel[8];
				ans[3231]<=tmp[3130]*kernel[0]+tmp[3131]*kernel[1]+tmp[3132]*kernel[2]+tmp[3230]*kernel[3]+tmp[3231]*kernel[4]+tmp[3232]*kernel[5]+tmp[3330]*kernel[6]+tmp[3331]*kernel[7]+tmp[3332]*kernel[8];
				ans[3232]<=tmp[3131]*kernel[0]+tmp[3132]*kernel[1]+tmp[3133]*kernel[2]+tmp[3231]*kernel[3]+tmp[3232]*kernel[4]+tmp[3233]*kernel[5]+tmp[3331]*kernel[6]+tmp[3332]*kernel[7]+tmp[3333]*kernel[8];
				ans[3233]<=tmp[3132]*kernel[0]+tmp[3133]*kernel[1]+tmp[3134]*kernel[2]+tmp[3232]*kernel[3]+tmp[3233]*kernel[4]+tmp[3234]*kernel[5]+tmp[3332]*kernel[6]+tmp[3333]*kernel[7]+tmp[3334]*kernel[8];
				ans[3234]<=tmp[3133]*kernel[0]+tmp[3134]*kernel[1]+tmp[3135]*kernel[2]+tmp[3233]*kernel[3]+tmp[3234]*kernel[4]+tmp[3235]*kernel[5]+tmp[3333]*kernel[6]+tmp[3334]*kernel[7]+tmp[3335]*kernel[8];
				ans[3235]<=tmp[3134]*kernel[0]+tmp[3135]*kernel[1]+tmp[3136]*kernel[2]+tmp[3234]*kernel[3]+tmp[3235]*kernel[4]+tmp[3236]*kernel[5]+tmp[3334]*kernel[6]+tmp[3335]*kernel[7]+tmp[3336]*kernel[8];
				ans[3236]<=tmp[3135]*kernel[0]+tmp[3136]*kernel[1]+tmp[3137]*kernel[2]+tmp[3235]*kernel[3]+tmp[3236]*kernel[4]+tmp[3237]*kernel[5]+tmp[3335]*kernel[6]+tmp[3336]*kernel[7]+tmp[3337]*kernel[8];
				ans[3237]<=tmp[3136]*kernel[0]+tmp[3137]*kernel[1]+tmp[3138]*kernel[2]+tmp[3236]*kernel[3]+tmp[3237]*kernel[4]+tmp[3238]*kernel[5]+tmp[3336]*kernel[6]+tmp[3337]*kernel[7]+tmp[3338]*kernel[8];
				ans[3238]<=tmp[3137]*kernel[0]+tmp[3138]*kernel[1]+tmp[3139]*kernel[2]+tmp[3237]*kernel[3]+tmp[3238]*kernel[4]+tmp[3239]*kernel[5]+tmp[3337]*kernel[6]+tmp[3338]*kernel[7]+tmp[3339]*kernel[8];
				ans[3239]<=tmp[3138]*kernel[0]+tmp[3139]*kernel[1]+tmp[3140]*kernel[2]+tmp[3238]*kernel[3]+tmp[3239]*kernel[4]+tmp[3240]*kernel[5]+tmp[3338]*kernel[6]+tmp[3339]*kernel[7]+tmp[3340]*kernel[8];
				ans[3240]<=tmp[3139]*kernel[0]+tmp[3140]*kernel[1]+tmp[3141]*kernel[2]+tmp[3239]*kernel[3]+tmp[3240]*kernel[4]+tmp[3241]*kernel[5]+tmp[3339]*kernel[6]+tmp[3340]*kernel[7]+tmp[3341]*kernel[8];
				ans[3241]<=tmp[3140]*kernel[0]+tmp[3141]*kernel[1]+tmp[3142]*kernel[2]+tmp[3240]*kernel[3]+tmp[3241]*kernel[4]+tmp[3242]*kernel[5]+tmp[3340]*kernel[6]+tmp[3341]*kernel[7]+tmp[3342]*kernel[8];
				ans[3242]<=tmp[3141]*kernel[0]+tmp[3142]*kernel[1]+tmp[3143]*kernel[2]+tmp[3241]*kernel[3]+tmp[3242]*kernel[4]+tmp[3243]*kernel[5]+tmp[3341]*kernel[6]+tmp[3342]*kernel[7]+tmp[3343]*kernel[8];
				ans[3243]<=tmp[3142]*kernel[0]+tmp[3143]*kernel[1]+tmp[3144]*kernel[2]+tmp[3242]*kernel[3]+tmp[3243]*kernel[4]+tmp[3244]*kernel[5]+tmp[3342]*kernel[6]+tmp[3343]*kernel[7]+tmp[3344]*kernel[8];
				ans[3244]<=tmp[3143]*kernel[0]+tmp[3144]*kernel[1]+tmp[3145]*kernel[2]+tmp[3243]*kernel[3]+tmp[3244]*kernel[4]+tmp[3245]*kernel[5]+tmp[3343]*kernel[6]+tmp[3344]*kernel[7]+tmp[3345]*kernel[8];
				ans[3245]<=tmp[3144]*kernel[0]+tmp[3145]*kernel[1]+tmp[3146]*kernel[2]+tmp[3244]*kernel[3]+tmp[3245]*kernel[4]+tmp[3246]*kernel[5]+tmp[3344]*kernel[6]+tmp[3345]*kernel[7]+tmp[3346]*kernel[8];
				ans[3246]<=tmp[3145]*kernel[0]+tmp[3146]*kernel[1]+tmp[3147]*kernel[2]+tmp[3245]*kernel[3]+tmp[3246]*kernel[4]+tmp[3247]*kernel[5]+tmp[3345]*kernel[6]+tmp[3346]*kernel[7]+tmp[3347]*kernel[8];
				ans[3247]<=tmp[3146]*kernel[0]+tmp[3147]*kernel[1]+tmp[3148]*kernel[2]+tmp[3246]*kernel[3]+tmp[3247]*kernel[4]+tmp[3248]*kernel[5]+tmp[3346]*kernel[6]+tmp[3347]*kernel[7]+tmp[3348]*kernel[8];
				ans[3248]<=tmp[3147]*kernel[0]+tmp[3148]*kernel[1]+tmp[3149]*kernel[2]+tmp[3247]*kernel[3]+tmp[3248]*kernel[4]+tmp[3249]*kernel[5]+tmp[3347]*kernel[6]+tmp[3348]*kernel[7]+tmp[3349]*kernel[8];
				ans[3249]<=tmp[3148]*kernel[0]+tmp[3149]*kernel[1]+tmp[3150]*kernel[2]+tmp[3248]*kernel[3]+tmp[3249]*kernel[4]+tmp[3250]*kernel[5]+tmp[3348]*kernel[6]+tmp[3349]*kernel[7]+tmp[3350]*kernel[8];
				ans[3250]<=tmp[3149]*kernel[0]+tmp[3150]*kernel[1]+tmp[3151]*kernel[2]+tmp[3249]*kernel[3]+tmp[3250]*kernel[4]+tmp[3251]*kernel[5]+tmp[3349]*kernel[6]+tmp[3350]*kernel[7]+tmp[3351]*kernel[8];
				ans[3251]<=tmp[3150]*kernel[0]+tmp[3151]*kernel[1]+tmp[3152]*kernel[2]+tmp[3250]*kernel[3]+tmp[3251]*kernel[4]+tmp[3252]*kernel[5]+tmp[3350]*kernel[6]+tmp[3351]*kernel[7]+tmp[3352]*kernel[8];
				ans[3252]<=tmp[3151]*kernel[0]+tmp[3152]*kernel[1]+tmp[3153]*kernel[2]+tmp[3251]*kernel[3]+tmp[3252]*kernel[4]+tmp[3253]*kernel[5]+tmp[3351]*kernel[6]+tmp[3352]*kernel[7]+tmp[3353]*kernel[8];
				ans[3253]<=tmp[3152]*kernel[0]+tmp[3153]*kernel[1]+tmp[3154]*kernel[2]+tmp[3252]*kernel[3]+tmp[3253]*kernel[4]+tmp[3254]*kernel[5]+tmp[3352]*kernel[6]+tmp[3353]*kernel[7]+tmp[3354]*kernel[8];
				ans[3254]<=tmp[3153]*kernel[0]+tmp[3154]*kernel[1]+tmp[3155]*kernel[2]+tmp[3253]*kernel[3]+tmp[3254]*kernel[4]+tmp[3255]*kernel[5]+tmp[3353]*kernel[6]+tmp[3354]*kernel[7]+tmp[3355]*kernel[8];
				ans[3255]<=tmp[3154]*kernel[0]+tmp[3155]*kernel[1]+tmp[3156]*kernel[2]+tmp[3254]*kernel[3]+tmp[3255]*kernel[4]+tmp[3256]*kernel[5]+tmp[3354]*kernel[6]+tmp[3355]*kernel[7]+tmp[3356]*kernel[8];
				ans[3256]<=tmp[3155]*kernel[0]+tmp[3156]*kernel[1]+tmp[3157]*kernel[2]+tmp[3255]*kernel[3]+tmp[3256]*kernel[4]+tmp[3257]*kernel[5]+tmp[3355]*kernel[6]+tmp[3356]*kernel[7]+tmp[3357]*kernel[8];
				ans[3257]<=tmp[3156]*kernel[0]+tmp[3157]*kernel[1]+tmp[3158]*kernel[2]+tmp[3256]*kernel[3]+tmp[3257]*kernel[4]+tmp[3258]*kernel[5]+tmp[3356]*kernel[6]+tmp[3357]*kernel[7]+tmp[3358]*kernel[8];
				ans[3258]<=tmp[3157]*kernel[0]+tmp[3158]*kernel[1]+tmp[3159]*kernel[2]+tmp[3257]*kernel[3]+tmp[3258]*kernel[4]+tmp[3259]*kernel[5]+tmp[3357]*kernel[6]+tmp[3358]*kernel[7]+tmp[3359]*kernel[8];
				ans[3259]<=tmp[3158]*kernel[0]+tmp[3159]*kernel[1]+tmp[3160]*kernel[2]+tmp[3258]*kernel[3]+tmp[3259]*kernel[4]+tmp[3260]*kernel[5]+tmp[3358]*kernel[6]+tmp[3359]*kernel[7]+tmp[3360]*kernel[8];
				ans[3260]<=tmp[3159]*kernel[0]+tmp[3160]*kernel[1]+tmp[3161]*kernel[2]+tmp[3259]*kernel[3]+tmp[3260]*kernel[4]+tmp[3261]*kernel[5]+tmp[3359]*kernel[6]+tmp[3360]*kernel[7]+tmp[3361]*kernel[8];
				ans[3261]<=tmp[3160]*kernel[0]+tmp[3161]*kernel[1]+tmp[3162]*kernel[2]+tmp[3260]*kernel[3]+tmp[3261]*kernel[4]+tmp[3262]*kernel[5]+tmp[3360]*kernel[6]+tmp[3361]*kernel[7]+tmp[3362]*kernel[8];
				ans[3262]<=tmp[3161]*kernel[0]+tmp[3162]*kernel[1]+tmp[3163]*kernel[2]+tmp[3261]*kernel[3]+tmp[3262]*kernel[4]+tmp[3263]*kernel[5]+tmp[3361]*kernel[6]+tmp[3362]*kernel[7]+tmp[3363]*kernel[8];
				ans[3263]<=tmp[3162]*kernel[0]+tmp[3163]*kernel[1]+tmp[3164]*kernel[2]+tmp[3262]*kernel[3]+tmp[3263]*kernel[4]+tmp[3264]*kernel[5]+tmp[3362]*kernel[6]+tmp[3363]*kernel[7]+tmp[3364]*kernel[8];
				ans[3264]<=tmp[3163]*kernel[0]+tmp[3164]*kernel[1]+tmp[3165]*kernel[2]+tmp[3263]*kernel[3]+tmp[3264]*kernel[4]+tmp[3265]*kernel[5]+tmp[3363]*kernel[6]+tmp[3364]*kernel[7]+tmp[3365]*kernel[8];
				ans[3265]<=tmp[3164]*kernel[0]+tmp[3165]*kernel[1]+tmp[3166]*kernel[2]+tmp[3264]*kernel[3]+tmp[3265]*kernel[4]+tmp[3266]*kernel[5]+tmp[3364]*kernel[6]+tmp[3365]*kernel[7]+tmp[3366]*kernel[8];
				ans[3266]<=tmp[3165]*kernel[0]+tmp[3166]*kernel[1]+tmp[3167]*kernel[2]+tmp[3265]*kernel[3]+tmp[3266]*kernel[4]+tmp[3267]*kernel[5]+tmp[3365]*kernel[6]+tmp[3366]*kernel[7]+tmp[3367]*kernel[8];
				ans[3267]<=tmp[3166]*kernel[0]+tmp[3167]*kernel[1]+tmp[3168]*kernel[2]+tmp[3266]*kernel[3]+tmp[3267]*kernel[4]+tmp[3268]*kernel[5]+tmp[3366]*kernel[6]+tmp[3367]*kernel[7]+tmp[3368]*kernel[8];
				ans[3268]<=tmp[3167]*kernel[0]+tmp[3168]*kernel[1]+tmp[3169]*kernel[2]+tmp[3267]*kernel[3]+tmp[3268]*kernel[4]+tmp[3269]*kernel[5]+tmp[3367]*kernel[6]+tmp[3368]*kernel[7]+tmp[3369]*kernel[8];
				ans[3269]<=tmp[3168]*kernel[0]+tmp[3169]*kernel[1]+tmp[3170]*kernel[2]+tmp[3268]*kernel[3]+tmp[3269]*kernel[4]+tmp[3270]*kernel[5]+tmp[3368]*kernel[6]+tmp[3369]*kernel[7]+tmp[3370]*kernel[8];
				ans[3270]<=tmp[3169]*kernel[0]+tmp[3170]*kernel[1]+tmp[3171]*kernel[2]+tmp[3269]*kernel[3]+tmp[3270]*kernel[4]+tmp[3271]*kernel[5]+tmp[3369]*kernel[6]+tmp[3370]*kernel[7]+tmp[3371]*kernel[8];
				ans[3271]<=tmp[3170]*kernel[0]+tmp[3171]*kernel[1]+tmp[3172]*kernel[2]+tmp[3270]*kernel[3]+tmp[3271]*kernel[4]+tmp[3272]*kernel[5]+tmp[3370]*kernel[6]+tmp[3371]*kernel[7]+tmp[3372]*kernel[8];
				ans[3272]<=tmp[3171]*kernel[0]+tmp[3172]*kernel[1]+tmp[3173]*kernel[2]+tmp[3271]*kernel[3]+tmp[3272]*kernel[4]+tmp[3273]*kernel[5]+tmp[3371]*kernel[6]+tmp[3372]*kernel[7]+tmp[3373]*kernel[8];
				ans[3273]<=tmp[3172]*kernel[0]+tmp[3173]*kernel[1]+tmp[3174]*kernel[2]+tmp[3272]*kernel[3]+tmp[3273]*kernel[4]+tmp[3274]*kernel[5]+tmp[3372]*kernel[6]+tmp[3373]*kernel[7]+tmp[3374]*kernel[8];
				ans[3274]<=tmp[3173]*kernel[0]+tmp[3174]*kernel[1]+tmp[3175]*kernel[2]+tmp[3273]*kernel[3]+tmp[3274]*kernel[4]+tmp[3275]*kernel[5]+tmp[3373]*kernel[6]+tmp[3374]*kernel[7]+tmp[3375]*kernel[8];
				ans[3275]<=tmp[3174]*kernel[0]+tmp[3175]*kernel[1]+tmp[3176]*kernel[2]+tmp[3274]*kernel[3]+tmp[3275]*kernel[4]+tmp[3276]*kernel[5]+tmp[3374]*kernel[6]+tmp[3375]*kernel[7]+tmp[3376]*kernel[8];
				ans[3276]<=tmp[3175]*kernel[0]+tmp[3176]*kernel[1]+tmp[3177]*kernel[2]+tmp[3275]*kernel[3]+tmp[3276]*kernel[4]+tmp[3277]*kernel[5]+tmp[3375]*kernel[6]+tmp[3376]*kernel[7]+tmp[3377]*kernel[8];
				ans[3277]<=tmp[3176]*kernel[0]+tmp[3177]*kernel[1]+tmp[3178]*kernel[2]+tmp[3276]*kernel[3]+tmp[3277]*kernel[4]+tmp[3278]*kernel[5]+tmp[3376]*kernel[6]+tmp[3377]*kernel[7]+tmp[3378]*kernel[8];
				ans[3278]<=tmp[3177]*kernel[0]+tmp[3178]*kernel[1]+tmp[3179]*kernel[2]+tmp[3277]*kernel[3]+tmp[3278]*kernel[4]+tmp[3279]*kernel[5]+tmp[3377]*kernel[6]+tmp[3378]*kernel[7]+tmp[3379]*kernel[8];
				ans[3279]<=tmp[3178]*kernel[0]+tmp[3179]*kernel[1]+tmp[3180]*kernel[2]+tmp[3278]*kernel[3]+tmp[3279]*kernel[4]+tmp[3280]*kernel[5]+tmp[3378]*kernel[6]+tmp[3379]*kernel[7]+tmp[3380]*kernel[8];
				ans[3280]<=tmp[3179]*kernel[0]+tmp[3180]*kernel[1]+tmp[3181]*kernel[2]+tmp[3279]*kernel[3]+tmp[3280]*kernel[4]+tmp[3281]*kernel[5]+tmp[3379]*kernel[6]+tmp[3380]*kernel[7]+tmp[3381]*kernel[8];
				ans[3281]<=tmp[3180]*kernel[0]+tmp[3181]*kernel[1]+tmp[3182]*kernel[2]+tmp[3280]*kernel[3]+tmp[3281]*kernel[4]+tmp[3282]*kernel[5]+tmp[3380]*kernel[6]+tmp[3381]*kernel[7]+tmp[3382]*kernel[8];
				ans[3282]<=tmp[3181]*kernel[0]+tmp[3182]*kernel[1]+tmp[3183]*kernel[2]+tmp[3281]*kernel[3]+tmp[3282]*kernel[4]+tmp[3283]*kernel[5]+tmp[3381]*kernel[6]+tmp[3382]*kernel[7]+tmp[3383]*kernel[8];
				ans[3283]<=tmp[3182]*kernel[0]+tmp[3183]*kernel[1]+tmp[3184]*kernel[2]+tmp[3282]*kernel[3]+tmp[3283]*kernel[4]+tmp[3284]*kernel[5]+tmp[3382]*kernel[6]+tmp[3383]*kernel[7]+tmp[3384]*kernel[8];
				ans[3284]<=tmp[3183]*kernel[0]+tmp[3184]*kernel[1]+tmp[3185]*kernel[2]+tmp[3283]*kernel[3]+tmp[3284]*kernel[4]+tmp[3285]*kernel[5]+tmp[3383]*kernel[6]+tmp[3384]*kernel[7]+tmp[3385]*kernel[8];
				ans[3285]<=tmp[3184]*kernel[0]+tmp[3185]*kernel[1]+tmp[3186]*kernel[2]+tmp[3284]*kernel[3]+tmp[3285]*kernel[4]+tmp[3286]*kernel[5]+tmp[3384]*kernel[6]+tmp[3385]*kernel[7]+tmp[3386]*kernel[8];
				ans[3286]<=tmp[3185]*kernel[0]+tmp[3186]*kernel[1]+tmp[3187]*kernel[2]+tmp[3285]*kernel[3]+tmp[3286]*kernel[4]+tmp[3287]*kernel[5]+tmp[3385]*kernel[6]+tmp[3386]*kernel[7]+tmp[3387]*kernel[8];
				ans[3287]<=tmp[3186]*kernel[0]+tmp[3187]*kernel[1]+tmp[3188]*kernel[2]+tmp[3286]*kernel[3]+tmp[3287]*kernel[4]+tmp[3288]*kernel[5]+tmp[3386]*kernel[6]+tmp[3387]*kernel[7]+tmp[3388]*kernel[8];
				ans[3288]<=tmp[3187]*kernel[0]+tmp[3188]*kernel[1]+tmp[3189]*kernel[2]+tmp[3287]*kernel[3]+tmp[3288]*kernel[4]+tmp[3289]*kernel[5]+tmp[3387]*kernel[6]+tmp[3388]*kernel[7]+tmp[3389]*kernel[8];
				ans[3289]<=tmp[3188]*kernel[0]+tmp[3189]*kernel[1]+tmp[3190]*kernel[2]+tmp[3288]*kernel[3]+tmp[3289]*kernel[4]+tmp[3290]*kernel[5]+tmp[3388]*kernel[6]+tmp[3389]*kernel[7]+tmp[3390]*kernel[8];
				ans[3290]<=tmp[3189]*kernel[0]+tmp[3190]*kernel[1]+tmp[3191]*kernel[2]+tmp[3289]*kernel[3]+tmp[3290]*kernel[4]+tmp[3291]*kernel[5]+tmp[3389]*kernel[6]+tmp[3390]*kernel[7]+tmp[3391]*kernel[8];
				ans[3291]<=tmp[3190]*kernel[0]+tmp[3191]*kernel[1]+tmp[3192]*kernel[2]+tmp[3290]*kernel[3]+tmp[3291]*kernel[4]+tmp[3292]*kernel[5]+tmp[3390]*kernel[6]+tmp[3391]*kernel[7]+tmp[3392]*kernel[8];
				ans[3292]<=tmp[3191]*kernel[0]+tmp[3192]*kernel[1]+tmp[3193]*kernel[2]+tmp[3291]*kernel[3]+tmp[3292]*kernel[4]+tmp[3293]*kernel[5]+tmp[3391]*kernel[6]+tmp[3392]*kernel[7]+tmp[3393]*kernel[8];
				ans[3293]<=tmp[3192]*kernel[0]+tmp[3193]*kernel[1]+tmp[3194]*kernel[2]+tmp[3292]*kernel[3]+tmp[3293]*kernel[4]+tmp[3294]*kernel[5]+tmp[3392]*kernel[6]+tmp[3393]*kernel[7]+tmp[3394]*kernel[8];
				ans[3294]<=tmp[3193]*kernel[0]+tmp[3194]*kernel[1]+tmp[3195]*kernel[2]+tmp[3293]*kernel[3]+tmp[3294]*kernel[4]+tmp[3295]*kernel[5]+tmp[3393]*kernel[6]+tmp[3394]*kernel[7]+tmp[3395]*kernel[8];
				ans[3295]<=tmp[3194]*kernel[0]+tmp[3195]*kernel[1]+tmp[3196]*kernel[2]+tmp[3294]*kernel[3]+tmp[3295]*kernel[4]+tmp[3296]*kernel[5]+tmp[3394]*kernel[6]+tmp[3395]*kernel[7]+tmp[3396]*kernel[8];
				ans[3296]<=tmp[3195]*kernel[0]+tmp[3196]*kernel[1]+tmp[3197]*kernel[2]+tmp[3295]*kernel[3]+tmp[3296]*kernel[4]+tmp[3297]*kernel[5]+tmp[3395]*kernel[6]+tmp[3396]*kernel[7]+tmp[3397]*kernel[8];
				ans[3297]<=tmp[3196]*kernel[0]+tmp[3197]*kernel[1]+tmp[3198]*kernel[2]+tmp[3296]*kernel[3]+tmp[3297]*kernel[4]+tmp[3298]*kernel[5]+tmp[3396]*kernel[6]+tmp[3397]*kernel[7]+tmp[3398]*kernel[8];
				ans[3298]<=tmp[3197]*kernel[0]+tmp[3198]*kernel[1]+tmp[3199]*kernel[2]+tmp[3297]*kernel[3]+tmp[3298]*kernel[4]+tmp[3299]*kernel[5]+tmp[3397]*kernel[6]+tmp[3398]*kernel[7]+tmp[3399]*kernel[8];
				ans[3299]<=tmp[3198]*kernel[0]+tmp[3199]*kernel[1]+tmp[3298]*kernel[3]+tmp[3299]*kernel[4]+tmp[3398]*kernel[6]+tmp[3399]*kernel[7];
				ans[3300]<=tmp[3200]*kernel[1]+tmp[3201]*kernel[2]+tmp[3300]*kernel[4]+tmp[3301]*kernel[5]+tmp[3400]*kernel[7]+tmp[3401]*kernel[8];
				ans[3301]<=tmp[3200]*kernel[0]+tmp[3201]*kernel[1]+tmp[3202]*kernel[2]+tmp[3300]*kernel[3]+tmp[3301]*kernel[4]+tmp[3302]*kernel[5]+tmp[3400]*kernel[6]+tmp[3401]*kernel[7]+tmp[3402]*kernel[8];
				ans[3302]<=tmp[3201]*kernel[0]+tmp[3202]*kernel[1]+tmp[3203]*kernel[2]+tmp[3301]*kernel[3]+tmp[3302]*kernel[4]+tmp[3303]*kernel[5]+tmp[3401]*kernel[6]+tmp[3402]*kernel[7]+tmp[3403]*kernel[8];
				ans[3303]<=tmp[3202]*kernel[0]+tmp[3203]*kernel[1]+tmp[3204]*kernel[2]+tmp[3302]*kernel[3]+tmp[3303]*kernel[4]+tmp[3304]*kernel[5]+tmp[3402]*kernel[6]+tmp[3403]*kernel[7]+tmp[3404]*kernel[8];
				ans[3304]<=tmp[3203]*kernel[0]+tmp[3204]*kernel[1]+tmp[3205]*kernel[2]+tmp[3303]*kernel[3]+tmp[3304]*kernel[4]+tmp[3305]*kernel[5]+tmp[3403]*kernel[6]+tmp[3404]*kernel[7]+tmp[3405]*kernel[8];
				ans[3305]<=tmp[3204]*kernel[0]+tmp[3205]*kernel[1]+tmp[3206]*kernel[2]+tmp[3304]*kernel[3]+tmp[3305]*kernel[4]+tmp[3306]*kernel[5]+tmp[3404]*kernel[6]+tmp[3405]*kernel[7]+tmp[3406]*kernel[8];
				ans[3306]<=tmp[3205]*kernel[0]+tmp[3206]*kernel[1]+tmp[3207]*kernel[2]+tmp[3305]*kernel[3]+tmp[3306]*kernel[4]+tmp[3307]*kernel[5]+tmp[3405]*kernel[6]+tmp[3406]*kernel[7]+tmp[3407]*kernel[8];
				ans[3307]<=tmp[3206]*kernel[0]+tmp[3207]*kernel[1]+tmp[3208]*kernel[2]+tmp[3306]*kernel[3]+tmp[3307]*kernel[4]+tmp[3308]*kernel[5]+tmp[3406]*kernel[6]+tmp[3407]*kernel[7]+tmp[3408]*kernel[8];
				ans[3308]<=tmp[3207]*kernel[0]+tmp[3208]*kernel[1]+tmp[3209]*kernel[2]+tmp[3307]*kernel[3]+tmp[3308]*kernel[4]+tmp[3309]*kernel[5]+tmp[3407]*kernel[6]+tmp[3408]*kernel[7]+tmp[3409]*kernel[8];
				ans[3309]<=tmp[3208]*kernel[0]+tmp[3209]*kernel[1]+tmp[3210]*kernel[2]+tmp[3308]*kernel[3]+tmp[3309]*kernel[4]+tmp[3310]*kernel[5]+tmp[3408]*kernel[6]+tmp[3409]*kernel[7]+tmp[3410]*kernel[8];
				ans[3310]<=tmp[3209]*kernel[0]+tmp[3210]*kernel[1]+tmp[3211]*kernel[2]+tmp[3309]*kernel[3]+tmp[3310]*kernel[4]+tmp[3311]*kernel[5]+tmp[3409]*kernel[6]+tmp[3410]*kernel[7]+tmp[3411]*kernel[8];
				ans[3311]<=tmp[3210]*kernel[0]+tmp[3211]*kernel[1]+tmp[3212]*kernel[2]+tmp[3310]*kernel[3]+tmp[3311]*kernel[4]+tmp[3312]*kernel[5]+tmp[3410]*kernel[6]+tmp[3411]*kernel[7]+tmp[3412]*kernel[8];
				ans[3312]<=tmp[3211]*kernel[0]+tmp[3212]*kernel[1]+tmp[3213]*kernel[2]+tmp[3311]*kernel[3]+tmp[3312]*kernel[4]+tmp[3313]*kernel[5]+tmp[3411]*kernel[6]+tmp[3412]*kernel[7]+tmp[3413]*kernel[8];
				ans[3313]<=tmp[3212]*kernel[0]+tmp[3213]*kernel[1]+tmp[3214]*kernel[2]+tmp[3312]*kernel[3]+tmp[3313]*kernel[4]+tmp[3314]*kernel[5]+tmp[3412]*kernel[6]+tmp[3413]*kernel[7]+tmp[3414]*kernel[8];
				ans[3314]<=tmp[3213]*kernel[0]+tmp[3214]*kernel[1]+tmp[3215]*kernel[2]+tmp[3313]*kernel[3]+tmp[3314]*kernel[4]+tmp[3315]*kernel[5]+tmp[3413]*kernel[6]+tmp[3414]*kernel[7]+tmp[3415]*kernel[8];
				ans[3315]<=tmp[3214]*kernel[0]+tmp[3215]*kernel[1]+tmp[3216]*kernel[2]+tmp[3314]*kernel[3]+tmp[3315]*kernel[4]+tmp[3316]*kernel[5]+tmp[3414]*kernel[6]+tmp[3415]*kernel[7]+tmp[3416]*kernel[8];
				ans[3316]<=tmp[3215]*kernel[0]+tmp[3216]*kernel[1]+tmp[3217]*kernel[2]+tmp[3315]*kernel[3]+tmp[3316]*kernel[4]+tmp[3317]*kernel[5]+tmp[3415]*kernel[6]+tmp[3416]*kernel[7]+tmp[3417]*kernel[8];
				ans[3317]<=tmp[3216]*kernel[0]+tmp[3217]*kernel[1]+tmp[3218]*kernel[2]+tmp[3316]*kernel[3]+tmp[3317]*kernel[4]+tmp[3318]*kernel[5]+tmp[3416]*kernel[6]+tmp[3417]*kernel[7]+tmp[3418]*kernel[8];
				ans[3318]<=tmp[3217]*kernel[0]+tmp[3218]*kernel[1]+tmp[3219]*kernel[2]+tmp[3317]*kernel[3]+tmp[3318]*kernel[4]+tmp[3319]*kernel[5]+tmp[3417]*kernel[6]+tmp[3418]*kernel[7]+tmp[3419]*kernel[8];
				ans[3319]<=tmp[3218]*kernel[0]+tmp[3219]*kernel[1]+tmp[3220]*kernel[2]+tmp[3318]*kernel[3]+tmp[3319]*kernel[4]+tmp[3320]*kernel[5]+tmp[3418]*kernel[6]+tmp[3419]*kernel[7]+tmp[3420]*kernel[8];
				ans[3320]<=tmp[3219]*kernel[0]+tmp[3220]*kernel[1]+tmp[3221]*kernel[2]+tmp[3319]*kernel[3]+tmp[3320]*kernel[4]+tmp[3321]*kernel[5]+tmp[3419]*kernel[6]+tmp[3420]*kernel[7]+tmp[3421]*kernel[8];
				ans[3321]<=tmp[3220]*kernel[0]+tmp[3221]*kernel[1]+tmp[3222]*kernel[2]+tmp[3320]*kernel[3]+tmp[3321]*kernel[4]+tmp[3322]*kernel[5]+tmp[3420]*kernel[6]+tmp[3421]*kernel[7]+tmp[3422]*kernel[8];
				ans[3322]<=tmp[3221]*kernel[0]+tmp[3222]*kernel[1]+tmp[3223]*kernel[2]+tmp[3321]*kernel[3]+tmp[3322]*kernel[4]+tmp[3323]*kernel[5]+tmp[3421]*kernel[6]+tmp[3422]*kernel[7]+tmp[3423]*kernel[8];
				ans[3323]<=tmp[3222]*kernel[0]+tmp[3223]*kernel[1]+tmp[3224]*kernel[2]+tmp[3322]*kernel[3]+tmp[3323]*kernel[4]+tmp[3324]*kernel[5]+tmp[3422]*kernel[6]+tmp[3423]*kernel[7]+tmp[3424]*kernel[8];
				ans[3324]<=tmp[3223]*kernel[0]+tmp[3224]*kernel[1]+tmp[3225]*kernel[2]+tmp[3323]*kernel[3]+tmp[3324]*kernel[4]+tmp[3325]*kernel[5]+tmp[3423]*kernel[6]+tmp[3424]*kernel[7]+tmp[3425]*kernel[8];
				ans[3325]<=tmp[3224]*kernel[0]+tmp[3225]*kernel[1]+tmp[3226]*kernel[2]+tmp[3324]*kernel[3]+tmp[3325]*kernel[4]+tmp[3326]*kernel[5]+tmp[3424]*kernel[6]+tmp[3425]*kernel[7]+tmp[3426]*kernel[8];
				ans[3326]<=tmp[3225]*kernel[0]+tmp[3226]*kernel[1]+tmp[3227]*kernel[2]+tmp[3325]*kernel[3]+tmp[3326]*kernel[4]+tmp[3327]*kernel[5]+tmp[3425]*kernel[6]+tmp[3426]*kernel[7]+tmp[3427]*kernel[8];
				ans[3327]<=tmp[3226]*kernel[0]+tmp[3227]*kernel[1]+tmp[3228]*kernel[2]+tmp[3326]*kernel[3]+tmp[3327]*kernel[4]+tmp[3328]*kernel[5]+tmp[3426]*kernel[6]+tmp[3427]*kernel[7]+tmp[3428]*kernel[8];
				ans[3328]<=tmp[3227]*kernel[0]+tmp[3228]*kernel[1]+tmp[3229]*kernel[2]+tmp[3327]*kernel[3]+tmp[3328]*kernel[4]+tmp[3329]*kernel[5]+tmp[3427]*kernel[6]+tmp[3428]*kernel[7]+tmp[3429]*kernel[8];
				ans[3329]<=tmp[3228]*kernel[0]+tmp[3229]*kernel[1]+tmp[3230]*kernel[2]+tmp[3328]*kernel[3]+tmp[3329]*kernel[4]+tmp[3330]*kernel[5]+tmp[3428]*kernel[6]+tmp[3429]*kernel[7]+tmp[3430]*kernel[8];
				ans[3330]<=tmp[3229]*kernel[0]+tmp[3230]*kernel[1]+tmp[3231]*kernel[2]+tmp[3329]*kernel[3]+tmp[3330]*kernel[4]+tmp[3331]*kernel[5]+tmp[3429]*kernel[6]+tmp[3430]*kernel[7]+tmp[3431]*kernel[8];
				ans[3331]<=tmp[3230]*kernel[0]+tmp[3231]*kernel[1]+tmp[3232]*kernel[2]+tmp[3330]*kernel[3]+tmp[3331]*kernel[4]+tmp[3332]*kernel[5]+tmp[3430]*kernel[6]+tmp[3431]*kernel[7]+tmp[3432]*kernel[8];
				ans[3332]<=tmp[3231]*kernel[0]+tmp[3232]*kernel[1]+tmp[3233]*kernel[2]+tmp[3331]*kernel[3]+tmp[3332]*kernel[4]+tmp[3333]*kernel[5]+tmp[3431]*kernel[6]+tmp[3432]*kernel[7]+tmp[3433]*kernel[8];
				ans[3333]<=tmp[3232]*kernel[0]+tmp[3233]*kernel[1]+tmp[3234]*kernel[2]+tmp[3332]*kernel[3]+tmp[3333]*kernel[4]+tmp[3334]*kernel[5]+tmp[3432]*kernel[6]+tmp[3433]*kernel[7]+tmp[3434]*kernel[8];
				ans[3334]<=tmp[3233]*kernel[0]+tmp[3234]*kernel[1]+tmp[3235]*kernel[2]+tmp[3333]*kernel[3]+tmp[3334]*kernel[4]+tmp[3335]*kernel[5]+tmp[3433]*kernel[6]+tmp[3434]*kernel[7]+tmp[3435]*kernel[8];
				ans[3335]<=tmp[3234]*kernel[0]+tmp[3235]*kernel[1]+tmp[3236]*kernel[2]+tmp[3334]*kernel[3]+tmp[3335]*kernel[4]+tmp[3336]*kernel[5]+tmp[3434]*kernel[6]+tmp[3435]*kernel[7]+tmp[3436]*kernel[8];
				ans[3336]<=tmp[3235]*kernel[0]+tmp[3236]*kernel[1]+tmp[3237]*kernel[2]+tmp[3335]*kernel[3]+tmp[3336]*kernel[4]+tmp[3337]*kernel[5]+tmp[3435]*kernel[6]+tmp[3436]*kernel[7]+tmp[3437]*kernel[8];
				ans[3337]<=tmp[3236]*kernel[0]+tmp[3237]*kernel[1]+tmp[3238]*kernel[2]+tmp[3336]*kernel[3]+tmp[3337]*kernel[4]+tmp[3338]*kernel[5]+tmp[3436]*kernel[6]+tmp[3437]*kernel[7]+tmp[3438]*kernel[8];
				ans[3338]<=tmp[3237]*kernel[0]+tmp[3238]*kernel[1]+tmp[3239]*kernel[2]+tmp[3337]*kernel[3]+tmp[3338]*kernel[4]+tmp[3339]*kernel[5]+tmp[3437]*kernel[6]+tmp[3438]*kernel[7]+tmp[3439]*kernel[8];
				ans[3339]<=tmp[3238]*kernel[0]+tmp[3239]*kernel[1]+tmp[3240]*kernel[2]+tmp[3338]*kernel[3]+tmp[3339]*kernel[4]+tmp[3340]*kernel[5]+tmp[3438]*kernel[6]+tmp[3439]*kernel[7]+tmp[3440]*kernel[8];
				ans[3340]<=tmp[3239]*kernel[0]+tmp[3240]*kernel[1]+tmp[3241]*kernel[2]+tmp[3339]*kernel[3]+tmp[3340]*kernel[4]+tmp[3341]*kernel[5]+tmp[3439]*kernel[6]+tmp[3440]*kernel[7]+tmp[3441]*kernel[8];
				ans[3341]<=tmp[3240]*kernel[0]+tmp[3241]*kernel[1]+tmp[3242]*kernel[2]+tmp[3340]*kernel[3]+tmp[3341]*kernel[4]+tmp[3342]*kernel[5]+tmp[3440]*kernel[6]+tmp[3441]*kernel[7]+tmp[3442]*kernel[8];
				ans[3342]<=tmp[3241]*kernel[0]+tmp[3242]*kernel[1]+tmp[3243]*kernel[2]+tmp[3341]*kernel[3]+tmp[3342]*kernel[4]+tmp[3343]*kernel[5]+tmp[3441]*kernel[6]+tmp[3442]*kernel[7]+tmp[3443]*kernel[8];
				ans[3343]<=tmp[3242]*kernel[0]+tmp[3243]*kernel[1]+tmp[3244]*kernel[2]+tmp[3342]*kernel[3]+tmp[3343]*kernel[4]+tmp[3344]*kernel[5]+tmp[3442]*kernel[6]+tmp[3443]*kernel[7]+tmp[3444]*kernel[8];
				ans[3344]<=tmp[3243]*kernel[0]+tmp[3244]*kernel[1]+tmp[3245]*kernel[2]+tmp[3343]*kernel[3]+tmp[3344]*kernel[4]+tmp[3345]*kernel[5]+tmp[3443]*kernel[6]+tmp[3444]*kernel[7]+tmp[3445]*kernel[8];
				ans[3345]<=tmp[3244]*kernel[0]+tmp[3245]*kernel[1]+tmp[3246]*kernel[2]+tmp[3344]*kernel[3]+tmp[3345]*kernel[4]+tmp[3346]*kernel[5]+tmp[3444]*kernel[6]+tmp[3445]*kernel[7]+tmp[3446]*kernel[8];
				ans[3346]<=tmp[3245]*kernel[0]+tmp[3246]*kernel[1]+tmp[3247]*kernel[2]+tmp[3345]*kernel[3]+tmp[3346]*kernel[4]+tmp[3347]*kernel[5]+tmp[3445]*kernel[6]+tmp[3446]*kernel[7]+tmp[3447]*kernel[8];
				ans[3347]<=tmp[3246]*kernel[0]+tmp[3247]*kernel[1]+tmp[3248]*kernel[2]+tmp[3346]*kernel[3]+tmp[3347]*kernel[4]+tmp[3348]*kernel[5]+tmp[3446]*kernel[6]+tmp[3447]*kernel[7]+tmp[3448]*kernel[8];
				ans[3348]<=tmp[3247]*kernel[0]+tmp[3248]*kernel[1]+tmp[3249]*kernel[2]+tmp[3347]*kernel[3]+tmp[3348]*kernel[4]+tmp[3349]*kernel[5]+tmp[3447]*kernel[6]+tmp[3448]*kernel[7]+tmp[3449]*kernel[8];
				ans[3349]<=tmp[3248]*kernel[0]+tmp[3249]*kernel[1]+tmp[3250]*kernel[2]+tmp[3348]*kernel[3]+tmp[3349]*kernel[4]+tmp[3350]*kernel[5]+tmp[3448]*kernel[6]+tmp[3449]*kernel[7]+tmp[3450]*kernel[8];
				ans[3350]<=tmp[3249]*kernel[0]+tmp[3250]*kernel[1]+tmp[3251]*kernel[2]+tmp[3349]*kernel[3]+tmp[3350]*kernel[4]+tmp[3351]*kernel[5]+tmp[3449]*kernel[6]+tmp[3450]*kernel[7]+tmp[3451]*kernel[8];
				ans[3351]<=tmp[3250]*kernel[0]+tmp[3251]*kernel[1]+tmp[3252]*kernel[2]+tmp[3350]*kernel[3]+tmp[3351]*kernel[4]+tmp[3352]*kernel[5]+tmp[3450]*kernel[6]+tmp[3451]*kernel[7]+tmp[3452]*kernel[8];
				ans[3352]<=tmp[3251]*kernel[0]+tmp[3252]*kernel[1]+tmp[3253]*kernel[2]+tmp[3351]*kernel[3]+tmp[3352]*kernel[4]+tmp[3353]*kernel[5]+tmp[3451]*kernel[6]+tmp[3452]*kernel[7]+tmp[3453]*kernel[8];
				ans[3353]<=tmp[3252]*kernel[0]+tmp[3253]*kernel[1]+tmp[3254]*kernel[2]+tmp[3352]*kernel[3]+tmp[3353]*kernel[4]+tmp[3354]*kernel[5]+tmp[3452]*kernel[6]+tmp[3453]*kernel[7]+tmp[3454]*kernel[8];
				ans[3354]<=tmp[3253]*kernel[0]+tmp[3254]*kernel[1]+tmp[3255]*kernel[2]+tmp[3353]*kernel[3]+tmp[3354]*kernel[4]+tmp[3355]*kernel[5]+tmp[3453]*kernel[6]+tmp[3454]*kernel[7]+tmp[3455]*kernel[8];
				ans[3355]<=tmp[3254]*kernel[0]+tmp[3255]*kernel[1]+tmp[3256]*kernel[2]+tmp[3354]*kernel[3]+tmp[3355]*kernel[4]+tmp[3356]*kernel[5]+tmp[3454]*kernel[6]+tmp[3455]*kernel[7]+tmp[3456]*kernel[8];
				ans[3356]<=tmp[3255]*kernel[0]+tmp[3256]*kernel[1]+tmp[3257]*kernel[2]+tmp[3355]*kernel[3]+tmp[3356]*kernel[4]+tmp[3357]*kernel[5]+tmp[3455]*kernel[6]+tmp[3456]*kernel[7]+tmp[3457]*kernel[8];
				ans[3357]<=tmp[3256]*kernel[0]+tmp[3257]*kernel[1]+tmp[3258]*kernel[2]+tmp[3356]*kernel[3]+tmp[3357]*kernel[4]+tmp[3358]*kernel[5]+tmp[3456]*kernel[6]+tmp[3457]*kernel[7]+tmp[3458]*kernel[8];
				ans[3358]<=tmp[3257]*kernel[0]+tmp[3258]*kernel[1]+tmp[3259]*kernel[2]+tmp[3357]*kernel[3]+tmp[3358]*kernel[4]+tmp[3359]*kernel[5]+tmp[3457]*kernel[6]+tmp[3458]*kernel[7]+tmp[3459]*kernel[8];
				ans[3359]<=tmp[3258]*kernel[0]+tmp[3259]*kernel[1]+tmp[3260]*kernel[2]+tmp[3358]*kernel[3]+tmp[3359]*kernel[4]+tmp[3360]*kernel[5]+tmp[3458]*kernel[6]+tmp[3459]*kernel[7]+tmp[3460]*kernel[8];
				ans[3360]<=tmp[3259]*kernel[0]+tmp[3260]*kernel[1]+tmp[3261]*kernel[2]+tmp[3359]*kernel[3]+tmp[3360]*kernel[4]+tmp[3361]*kernel[5]+tmp[3459]*kernel[6]+tmp[3460]*kernel[7]+tmp[3461]*kernel[8];
				ans[3361]<=tmp[3260]*kernel[0]+tmp[3261]*kernel[1]+tmp[3262]*kernel[2]+tmp[3360]*kernel[3]+tmp[3361]*kernel[4]+tmp[3362]*kernel[5]+tmp[3460]*kernel[6]+tmp[3461]*kernel[7]+tmp[3462]*kernel[8];
				ans[3362]<=tmp[3261]*kernel[0]+tmp[3262]*kernel[1]+tmp[3263]*kernel[2]+tmp[3361]*kernel[3]+tmp[3362]*kernel[4]+tmp[3363]*kernel[5]+tmp[3461]*kernel[6]+tmp[3462]*kernel[7]+tmp[3463]*kernel[8];
				ans[3363]<=tmp[3262]*kernel[0]+tmp[3263]*kernel[1]+tmp[3264]*kernel[2]+tmp[3362]*kernel[3]+tmp[3363]*kernel[4]+tmp[3364]*kernel[5]+tmp[3462]*kernel[6]+tmp[3463]*kernel[7]+tmp[3464]*kernel[8];
				ans[3364]<=tmp[3263]*kernel[0]+tmp[3264]*kernel[1]+tmp[3265]*kernel[2]+tmp[3363]*kernel[3]+tmp[3364]*kernel[4]+tmp[3365]*kernel[5]+tmp[3463]*kernel[6]+tmp[3464]*kernel[7]+tmp[3465]*kernel[8];
				ans[3365]<=tmp[3264]*kernel[0]+tmp[3265]*kernel[1]+tmp[3266]*kernel[2]+tmp[3364]*kernel[3]+tmp[3365]*kernel[4]+tmp[3366]*kernel[5]+tmp[3464]*kernel[6]+tmp[3465]*kernel[7]+tmp[3466]*kernel[8];
				ans[3366]<=tmp[3265]*kernel[0]+tmp[3266]*kernel[1]+tmp[3267]*kernel[2]+tmp[3365]*kernel[3]+tmp[3366]*kernel[4]+tmp[3367]*kernel[5]+tmp[3465]*kernel[6]+tmp[3466]*kernel[7]+tmp[3467]*kernel[8];
				ans[3367]<=tmp[3266]*kernel[0]+tmp[3267]*kernel[1]+tmp[3268]*kernel[2]+tmp[3366]*kernel[3]+tmp[3367]*kernel[4]+tmp[3368]*kernel[5]+tmp[3466]*kernel[6]+tmp[3467]*kernel[7]+tmp[3468]*kernel[8];
				ans[3368]<=tmp[3267]*kernel[0]+tmp[3268]*kernel[1]+tmp[3269]*kernel[2]+tmp[3367]*kernel[3]+tmp[3368]*kernel[4]+tmp[3369]*kernel[5]+tmp[3467]*kernel[6]+tmp[3468]*kernel[7]+tmp[3469]*kernel[8];
				ans[3369]<=tmp[3268]*kernel[0]+tmp[3269]*kernel[1]+tmp[3270]*kernel[2]+tmp[3368]*kernel[3]+tmp[3369]*kernel[4]+tmp[3370]*kernel[5]+tmp[3468]*kernel[6]+tmp[3469]*kernel[7]+tmp[3470]*kernel[8];
				ans[3370]<=tmp[3269]*kernel[0]+tmp[3270]*kernel[1]+tmp[3271]*kernel[2]+tmp[3369]*kernel[3]+tmp[3370]*kernel[4]+tmp[3371]*kernel[5]+tmp[3469]*kernel[6]+tmp[3470]*kernel[7]+tmp[3471]*kernel[8];
				ans[3371]<=tmp[3270]*kernel[0]+tmp[3271]*kernel[1]+tmp[3272]*kernel[2]+tmp[3370]*kernel[3]+tmp[3371]*kernel[4]+tmp[3372]*kernel[5]+tmp[3470]*kernel[6]+tmp[3471]*kernel[7]+tmp[3472]*kernel[8];
				ans[3372]<=tmp[3271]*kernel[0]+tmp[3272]*kernel[1]+tmp[3273]*kernel[2]+tmp[3371]*kernel[3]+tmp[3372]*kernel[4]+tmp[3373]*kernel[5]+tmp[3471]*kernel[6]+tmp[3472]*kernel[7]+tmp[3473]*kernel[8];
				ans[3373]<=tmp[3272]*kernel[0]+tmp[3273]*kernel[1]+tmp[3274]*kernel[2]+tmp[3372]*kernel[3]+tmp[3373]*kernel[4]+tmp[3374]*kernel[5]+tmp[3472]*kernel[6]+tmp[3473]*kernel[7]+tmp[3474]*kernel[8];
				ans[3374]<=tmp[3273]*kernel[0]+tmp[3274]*kernel[1]+tmp[3275]*kernel[2]+tmp[3373]*kernel[3]+tmp[3374]*kernel[4]+tmp[3375]*kernel[5]+tmp[3473]*kernel[6]+tmp[3474]*kernel[7]+tmp[3475]*kernel[8];
				ans[3375]<=tmp[3274]*kernel[0]+tmp[3275]*kernel[1]+tmp[3276]*kernel[2]+tmp[3374]*kernel[3]+tmp[3375]*kernel[4]+tmp[3376]*kernel[5]+tmp[3474]*kernel[6]+tmp[3475]*kernel[7]+tmp[3476]*kernel[8];
				ans[3376]<=tmp[3275]*kernel[0]+tmp[3276]*kernel[1]+tmp[3277]*kernel[2]+tmp[3375]*kernel[3]+tmp[3376]*kernel[4]+tmp[3377]*kernel[5]+tmp[3475]*kernel[6]+tmp[3476]*kernel[7]+tmp[3477]*kernel[8];
				ans[3377]<=tmp[3276]*kernel[0]+tmp[3277]*kernel[1]+tmp[3278]*kernel[2]+tmp[3376]*kernel[3]+tmp[3377]*kernel[4]+tmp[3378]*kernel[5]+tmp[3476]*kernel[6]+tmp[3477]*kernel[7]+tmp[3478]*kernel[8];
				ans[3378]<=tmp[3277]*kernel[0]+tmp[3278]*kernel[1]+tmp[3279]*kernel[2]+tmp[3377]*kernel[3]+tmp[3378]*kernel[4]+tmp[3379]*kernel[5]+tmp[3477]*kernel[6]+tmp[3478]*kernel[7]+tmp[3479]*kernel[8];
				ans[3379]<=tmp[3278]*kernel[0]+tmp[3279]*kernel[1]+tmp[3280]*kernel[2]+tmp[3378]*kernel[3]+tmp[3379]*kernel[4]+tmp[3380]*kernel[5]+tmp[3478]*kernel[6]+tmp[3479]*kernel[7]+tmp[3480]*kernel[8];
				ans[3380]<=tmp[3279]*kernel[0]+tmp[3280]*kernel[1]+tmp[3281]*kernel[2]+tmp[3379]*kernel[3]+tmp[3380]*kernel[4]+tmp[3381]*kernel[5]+tmp[3479]*kernel[6]+tmp[3480]*kernel[7]+tmp[3481]*kernel[8];
				ans[3381]<=tmp[3280]*kernel[0]+tmp[3281]*kernel[1]+tmp[3282]*kernel[2]+tmp[3380]*kernel[3]+tmp[3381]*kernel[4]+tmp[3382]*kernel[5]+tmp[3480]*kernel[6]+tmp[3481]*kernel[7]+tmp[3482]*kernel[8];
				ans[3382]<=tmp[3281]*kernel[0]+tmp[3282]*kernel[1]+tmp[3283]*kernel[2]+tmp[3381]*kernel[3]+tmp[3382]*kernel[4]+tmp[3383]*kernel[5]+tmp[3481]*kernel[6]+tmp[3482]*kernel[7]+tmp[3483]*kernel[8];
				ans[3383]<=tmp[3282]*kernel[0]+tmp[3283]*kernel[1]+tmp[3284]*kernel[2]+tmp[3382]*kernel[3]+tmp[3383]*kernel[4]+tmp[3384]*kernel[5]+tmp[3482]*kernel[6]+tmp[3483]*kernel[7]+tmp[3484]*kernel[8];
				ans[3384]<=tmp[3283]*kernel[0]+tmp[3284]*kernel[1]+tmp[3285]*kernel[2]+tmp[3383]*kernel[3]+tmp[3384]*kernel[4]+tmp[3385]*kernel[5]+tmp[3483]*kernel[6]+tmp[3484]*kernel[7]+tmp[3485]*kernel[8];
				ans[3385]<=tmp[3284]*kernel[0]+tmp[3285]*kernel[1]+tmp[3286]*kernel[2]+tmp[3384]*kernel[3]+tmp[3385]*kernel[4]+tmp[3386]*kernel[5]+tmp[3484]*kernel[6]+tmp[3485]*kernel[7]+tmp[3486]*kernel[8];
				ans[3386]<=tmp[3285]*kernel[0]+tmp[3286]*kernel[1]+tmp[3287]*kernel[2]+tmp[3385]*kernel[3]+tmp[3386]*kernel[4]+tmp[3387]*kernel[5]+tmp[3485]*kernel[6]+tmp[3486]*kernel[7]+tmp[3487]*kernel[8];
				ans[3387]<=tmp[3286]*kernel[0]+tmp[3287]*kernel[1]+tmp[3288]*kernel[2]+tmp[3386]*kernel[3]+tmp[3387]*kernel[4]+tmp[3388]*kernel[5]+tmp[3486]*kernel[6]+tmp[3487]*kernel[7]+tmp[3488]*kernel[8];
				ans[3388]<=tmp[3287]*kernel[0]+tmp[3288]*kernel[1]+tmp[3289]*kernel[2]+tmp[3387]*kernel[3]+tmp[3388]*kernel[4]+tmp[3389]*kernel[5]+tmp[3487]*kernel[6]+tmp[3488]*kernel[7]+tmp[3489]*kernel[8];
				ans[3389]<=tmp[3288]*kernel[0]+tmp[3289]*kernel[1]+tmp[3290]*kernel[2]+tmp[3388]*kernel[3]+tmp[3389]*kernel[4]+tmp[3390]*kernel[5]+tmp[3488]*kernel[6]+tmp[3489]*kernel[7]+tmp[3490]*kernel[8];
				ans[3390]<=tmp[3289]*kernel[0]+tmp[3290]*kernel[1]+tmp[3291]*kernel[2]+tmp[3389]*kernel[3]+tmp[3390]*kernel[4]+tmp[3391]*kernel[5]+tmp[3489]*kernel[6]+tmp[3490]*kernel[7]+tmp[3491]*kernel[8];
				ans[3391]<=tmp[3290]*kernel[0]+tmp[3291]*kernel[1]+tmp[3292]*kernel[2]+tmp[3390]*kernel[3]+tmp[3391]*kernel[4]+tmp[3392]*kernel[5]+tmp[3490]*kernel[6]+tmp[3491]*kernel[7]+tmp[3492]*kernel[8];
				ans[3392]<=tmp[3291]*kernel[0]+tmp[3292]*kernel[1]+tmp[3293]*kernel[2]+tmp[3391]*kernel[3]+tmp[3392]*kernel[4]+tmp[3393]*kernel[5]+tmp[3491]*kernel[6]+tmp[3492]*kernel[7]+tmp[3493]*kernel[8];
				ans[3393]<=tmp[3292]*kernel[0]+tmp[3293]*kernel[1]+tmp[3294]*kernel[2]+tmp[3392]*kernel[3]+tmp[3393]*kernel[4]+tmp[3394]*kernel[5]+tmp[3492]*kernel[6]+tmp[3493]*kernel[7]+tmp[3494]*kernel[8];
				ans[3394]<=tmp[3293]*kernel[0]+tmp[3294]*kernel[1]+tmp[3295]*kernel[2]+tmp[3393]*kernel[3]+tmp[3394]*kernel[4]+tmp[3395]*kernel[5]+tmp[3493]*kernel[6]+tmp[3494]*kernel[7]+tmp[3495]*kernel[8];
				ans[3395]<=tmp[3294]*kernel[0]+tmp[3295]*kernel[1]+tmp[3296]*kernel[2]+tmp[3394]*kernel[3]+tmp[3395]*kernel[4]+tmp[3396]*kernel[5]+tmp[3494]*kernel[6]+tmp[3495]*kernel[7]+tmp[3496]*kernel[8];
				ans[3396]<=tmp[3295]*kernel[0]+tmp[3296]*kernel[1]+tmp[3297]*kernel[2]+tmp[3395]*kernel[3]+tmp[3396]*kernel[4]+tmp[3397]*kernel[5]+tmp[3495]*kernel[6]+tmp[3496]*kernel[7]+tmp[3497]*kernel[8];
				ans[3397]<=tmp[3296]*kernel[0]+tmp[3297]*kernel[1]+tmp[3298]*kernel[2]+tmp[3396]*kernel[3]+tmp[3397]*kernel[4]+tmp[3398]*kernel[5]+tmp[3496]*kernel[6]+tmp[3497]*kernel[7]+tmp[3498]*kernel[8];
				ans[3398]<=tmp[3297]*kernel[0]+tmp[3298]*kernel[1]+tmp[3299]*kernel[2]+tmp[3397]*kernel[3]+tmp[3398]*kernel[4]+tmp[3399]*kernel[5]+tmp[3497]*kernel[6]+tmp[3498]*kernel[7]+tmp[3499]*kernel[8];
				ans[3399]<=tmp[3298]*kernel[0]+tmp[3299]*kernel[1]+tmp[3398]*kernel[3]+tmp[3399]*kernel[4]+tmp[3498]*kernel[6]+tmp[3499]*kernel[7];
				ans[3400]<=tmp[3300]*kernel[1]+tmp[3301]*kernel[2]+tmp[3400]*kernel[4]+tmp[3401]*kernel[5]+tmp[3500]*kernel[7]+tmp[3501]*kernel[8];
				ans[3401]<=tmp[3300]*kernel[0]+tmp[3301]*kernel[1]+tmp[3302]*kernel[2]+tmp[3400]*kernel[3]+tmp[3401]*kernel[4]+tmp[3402]*kernel[5]+tmp[3500]*kernel[6]+tmp[3501]*kernel[7]+tmp[3502]*kernel[8];
				ans[3402]<=tmp[3301]*kernel[0]+tmp[3302]*kernel[1]+tmp[3303]*kernel[2]+tmp[3401]*kernel[3]+tmp[3402]*kernel[4]+tmp[3403]*kernel[5]+tmp[3501]*kernel[6]+tmp[3502]*kernel[7]+tmp[3503]*kernel[8];
				ans[3403]<=tmp[3302]*kernel[0]+tmp[3303]*kernel[1]+tmp[3304]*kernel[2]+tmp[3402]*kernel[3]+tmp[3403]*kernel[4]+tmp[3404]*kernel[5]+tmp[3502]*kernel[6]+tmp[3503]*kernel[7]+tmp[3504]*kernel[8];
				ans[3404]<=tmp[3303]*kernel[0]+tmp[3304]*kernel[1]+tmp[3305]*kernel[2]+tmp[3403]*kernel[3]+tmp[3404]*kernel[4]+tmp[3405]*kernel[5]+tmp[3503]*kernel[6]+tmp[3504]*kernel[7]+tmp[3505]*kernel[8];
				ans[3405]<=tmp[3304]*kernel[0]+tmp[3305]*kernel[1]+tmp[3306]*kernel[2]+tmp[3404]*kernel[3]+tmp[3405]*kernel[4]+tmp[3406]*kernel[5]+tmp[3504]*kernel[6]+tmp[3505]*kernel[7]+tmp[3506]*kernel[8];
				ans[3406]<=tmp[3305]*kernel[0]+tmp[3306]*kernel[1]+tmp[3307]*kernel[2]+tmp[3405]*kernel[3]+tmp[3406]*kernel[4]+tmp[3407]*kernel[5]+tmp[3505]*kernel[6]+tmp[3506]*kernel[7]+tmp[3507]*kernel[8];
				ans[3407]<=tmp[3306]*kernel[0]+tmp[3307]*kernel[1]+tmp[3308]*kernel[2]+tmp[3406]*kernel[3]+tmp[3407]*kernel[4]+tmp[3408]*kernel[5]+tmp[3506]*kernel[6]+tmp[3507]*kernel[7]+tmp[3508]*kernel[8];
				ans[3408]<=tmp[3307]*kernel[0]+tmp[3308]*kernel[1]+tmp[3309]*kernel[2]+tmp[3407]*kernel[3]+tmp[3408]*kernel[4]+tmp[3409]*kernel[5]+tmp[3507]*kernel[6]+tmp[3508]*kernel[7]+tmp[3509]*kernel[8];
				ans[3409]<=tmp[3308]*kernel[0]+tmp[3309]*kernel[1]+tmp[3310]*kernel[2]+tmp[3408]*kernel[3]+tmp[3409]*kernel[4]+tmp[3410]*kernel[5]+tmp[3508]*kernel[6]+tmp[3509]*kernel[7]+tmp[3510]*kernel[8];
				ans[3410]<=tmp[3309]*kernel[0]+tmp[3310]*kernel[1]+tmp[3311]*kernel[2]+tmp[3409]*kernel[3]+tmp[3410]*kernel[4]+tmp[3411]*kernel[5]+tmp[3509]*kernel[6]+tmp[3510]*kernel[7]+tmp[3511]*kernel[8];
				ans[3411]<=tmp[3310]*kernel[0]+tmp[3311]*kernel[1]+tmp[3312]*kernel[2]+tmp[3410]*kernel[3]+tmp[3411]*kernel[4]+tmp[3412]*kernel[5]+tmp[3510]*kernel[6]+tmp[3511]*kernel[7]+tmp[3512]*kernel[8];
				ans[3412]<=tmp[3311]*kernel[0]+tmp[3312]*kernel[1]+tmp[3313]*kernel[2]+tmp[3411]*kernel[3]+tmp[3412]*kernel[4]+tmp[3413]*kernel[5]+tmp[3511]*kernel[6]+tmp[3512]*kernel[7]+tmp[3513]*kernel[8];
				ans[3413]<=tmp[3312]*kernel[0]+tmp[3313]*kernel[1]+tmp[3314]*kernel[2]+tmp[3412]*kernel[3]+tmp[3413]*kernel[4]+tmp[3414]*kernel[5]+tmp[3512]*kernel[6]+tmp[3513]*kernel[7]+tmp[3514]*kernel[8];
				ans[3414]<=tmp[3313]*kernel[0]+tmp[3314]*kernel[1]+tmp[3315]*kernel[2]+tmp[3413]*kernel[3]+tmp[3414]*kernel[4]+tmp[3415]*kernel[5]+tmp[3513]*kernel[6]+tmp[3514]*kernel[7]+tmp[3515]*kernel[8];
				ans[3415]<=tmp[3314]*kernel[0]+tmp[3315]*kernel[1]+tmp[3316]*kernel[2]+tmp[3414]*kernel[3]+tmp[3415]*kernel[4]+tmp[3416]*kernel[5]+tmp[3514]*kernel[6]+tmp[3515]*kernel[7]+tmp[3516]*kernel[8];
				ans[3416]<=tmp[3315]*kernel[0]+tmp[3316]*kernel[1]+tmp[3317]*kernel[2]+tmp[3415]*kernel[3]+tmp[3416]*kernel[4]+tmp[3417]*kernel[5]+tmp[3515]*kernel[6]+tmp[3516]*kernel[7]+tmp[3517]*kernel[8];
				ans[3417]<=tmp[3316]*kernel[0]+tmp[3317]*kernel[1]+tmp[3318]*kernel[2]+tmp[3416]*kernel[3]+tmp[3417]*kernel[4]+tmp[3418]*kernel[5]+tmp[3516]*kernel[6]+tmp[3517]*kernel[7]+tmp[3518]*kernel[8];
				ans[3418]<=tmp[3317]*kernel[0]+tmp[3318]*kernel[1]+tmp[3319]*kernel[2]+tmp[3417]*kernel[3]+tmp[3418]*kernel[4]+tmp[3419]*kernel[5]+tmp[3517]*kernel[6]+tmp[3518]*kernel[7]+tmp[3519]*kernel[8];
				ans[3419]<=tmp[3318]*kernel[0]+tmp[3319]*kernel[1]+tmp[3320]*kernel[2]+tmp[3418]*kernel[3]+tmp[3419]*kernel[4]+tmp[3420]*kernel[5]+tmp[3518]*kernel[6]+tmp[3519]*kernel[7]+tmp[3520]*kernel[8];
				ans[3420]<=tmp[3319]*kernel[0]+tmp[3320]*kernel[1]+tmp[3321]*kernel[2]+tmp[3419]*kernel[3]+tmp[3420]*kernel[4]+tmp[3421]*kernel[5]+tmp[3519]*kernel[6]+tmp[3520]*kernel[7]+tmp[3521]*kernel[8];
				ans[3421]<=tmp[3320]*kernel[0]+tmp[3321]*kernel[1]+tmp[3322]*kernel[2]+tmp[3420]*kernel[3]+tmp[3421]*kernel[4]+tmp[3422]*kernel[5]+tmp[3520]*kernel[6]+tmp[3521]*kernel[7]+tmp[3522]*kernel[8];
				ans[3422]<=tmp[3321]*kernel[0]+tmp[3322]*kernel[1]+tmp[3323]*kernel[2]+tmp[3421]*kernel[3]+tmp[3422]*kernel[4]+tmp[3423]*kernel[5]+tmp[3521]*kernel[6]+tmp[3522]*kernel[7]+tmp[3523]*kernel[8];
				ans[3423]<=tmp[3322]*kernel[0]+tmp[3323]*kernel[1]+tmp[3324]*kernel[2]+tmp[3422]*kernel[3]+tmp[3423]*kernel[4]+tmp[3424]*kernel[5]+tmp[3522]*kernel[6]+tmp[3523]*kernel[7]+tmp[3524]*kernel[8];
				ans[3424]<=tmp[3323]*kernel[0]+tmp[3324]*kernel[1]+tmp[3325]*kernel[2]+tmp[3423]*kernel[3]+tmp[3424]*kernel[4]+tmp[3425]*kernel[5]+tmp[3523]*kernel[6]+tmp[3524]*kernel[7]+tmp[3525]*kernel[8];
				ans[3425]<=tmp[3324]*kernel[0]+tmp[3325]*kernel[1]+tmp[3326]*kernel[2]+tmp[3424]*kernel[3]+tmp[3425]*kernel[4]+tmp[3426]*kernel[5]+tmp[3524]*kernel[6]+tmp[3525]*kernel[7]+tmp[3526]*kernel[8];
				ans[3426]<=tmp[3325]*kernel[0]+tmp[3326]*kernel[1]+tmp[3327]*kernel[2]+tmp[3425]*kernel[3]+tmp[3426]*kernel[4]+tmp[3427]*kernel[5]+tmp[3525]*kernel[6]+tmp[3526]*kernel[7]+tmp[3527]*kernel[8];
				ans[3427]<=tmp[3326]*kernel[0]+tmp[3327]*kernel[1]+tmp[3328]*kernel[2]+tmp[3426]*kernel[3]+tmp[3427]*kernel[4]+tmp[3428]*kernel[5]+tmp[3526]*kernel[6]+tmp[3527]*kernel[7]+tmp[3528]*kernel[8];
				ans[3428]<=tmp[3327]*kernel[0]+tmp[3328]*kernel[1]+tmp[3329]*kernel[2]+tmp[3427]*kernel[3]+tmp[3428]*kernel[4]+tmp[3429]*kernel[5]+tmp[3527]*kernel[6]+tmp[3528]*kernel[7]+tmp[3529]*kernel[8];
				ans[3429]<=tmp[3328]*kernel[0]+tmp[3329]*kernel[1]+tmp[3330]*kernel[2]+tmp[3428]*kernel[3]+tmp[3429]*kernel[4]+tmp[3430]*kernel[5]+tmp[3528]*kernel[6]+tmp[3529]*kernel[7]+tmp[3530]*kernel[8];
				ans[3430]<=tmp[3329]*kernel[0]+tmp[3330]*kernel[1]+tmp[3331]*kernel[2]+tmp[3429]*kernel[3]+tmp[3430]*kernel[4]+tmp[3431]*kernel[5]+tmp[3529]*kernel[6]+tmp[3530]*kernel[7]+tmp[3531]*kernel[8];
				ans[3431]<=tmp[3330]*kernel[0]+tmp[3331]*kernel[1]+tmp[3332]*kernel[2]+tmp[3430]*kernel[3]+tmp[3431]*kernel[4]+tmp[3432]*kernel[5]+tmp[3530]*kernel[6]+tmp[3531]*kernel[7]+tmp[3532]*kernel[8];
				ans[3432]<=tmp[3331]*kernel[0]+tmp[3332]*kernel[1]+tmp[3333]*kernel[2]+tmp[3431]*kernel[3]+tmp[3432]*kernel[4]+tmp[3433]*kernel[5]+tmp[3531]*kernel[6]+tmp[3532]*kernel[7]+tmp[3533]*kernel[8];
				ans[3433]<=tmp[3332]*kernel[0]+tmp[3333]*kernel[1]+tmp[3334]*kernel[2]+tmp[3432]*kernel[3]+tmp[3433]*kernel[4]+tmp[3434]*kernel[5]+tmp[3532]*kernel[6]+tmp[3533]*kernel[7]+tmp[3534]*kernel[8];
				ans[3434]<=tmp[3333]*kernel[0]+tmp[3334]*kernel[1]+tmp[3335]*kernel[2]+tmp[3433]*kernel[3]+tmp[3434]*kernel[4]+tmp[3435]*kernel[5]+tmp[3533]*kernel[6]+tmp[3534]*kernel[7]+tmp[3535]*kernel[8];
				ans[3435]<=tmp[3334]*kernel[0]+tmp[3335]*kernel[1]+tmp[3336]*kernel[2]+tmp[3434]*kernel[3]+tmp[3435]*kernel[4]+tmp[3436]*kernel[5]+tmp[3534]*kernel[6]+tmp[3535]*kernel[7]+tmp[3536]*kernel[8];
				ans[3436]<=tmp[3335]*kernel[0]+tmp[3336]*kernel[1]+tmp[3337]*kernel[2]+tmp[3435]*kernel[3]+tmp[3436]*kernel[4]+tmp[3437]*kernel[5]+tmp[3535]*kernel[6]+tmp[3536]*kernel[7]+tmp[3537]*kernel[8];
				ans[3437]<=tmp[3336]*kernel[0]+tmp[3337]*kernel[1]+tmp[3338]*kernel[2]+tmp[3436]*kernel[3]+tmp[3437]*kernel[4]+tmp[3438]*kernel[5]+tmp[3536]*kernel[6]+tmp[3537]*kernel[7]+tmp[3538]*kernel[8];
				ans[3438]<=tmp[3337]*kernel[0]+tmp[3338]*kernel[1]+tmp[3339]*kernel[2]+tmp[3437]*kernel[3]+tmp[3438]*kernel[4]+tmp[3439]*kernel[5]+tmp[3537]*kernel[6]+tmp[3538]*kernel[7]+tmp[3539]*kernel[8];
				ans[3439]<=tmp[3338]*kernel[0]+tmp[3339]*kernel[1]+tmp[3340]*kernel[2]+tmp[3438]*kernel[3]+tmp[3439]*kernel[4]+tmp[3440]*kernel[5]+tmp[3538]*kernel[6]+tmp[3539]*kernel[7]+tmp[3540]*kernel[8];
				ans[3440]<=tmp[3339]*kernel[0]+tmp[3340]*kernel[1]+tmp[3341]*kernel[2]+tmp[3439]*kernel[3]+tmp[3440]*kernel[4]+tmp[3441]*kernel[5]+tmp[3539]*kernel[6]+tmp[3540]*kernel[7]+tmp[3541]*kernel[8];
				ans[3441]<=tmp[3340]*kernel[0]+tmp[3341]*kernel[1]+tmp[3342]*kernel[2]+tmp[3440]*kernel[3]+tmp[3441]*kernel[4]+tmp[3442]*kernel[5]+tmp[3540]*kernel[6]+tmp[3541]*kernel[7]+tmp[3542]*kernel[8];
				ans[3442]<=tmp[3341]*kernel[0]+tmp[3342]*kernel[1]+tmp[3343]*kernel[2]+tmp[3441]*kernel[3]+tmp[3442]*kernel[4]+tmp[3443]*kernel[5]+tmp[3541]*kernel[6]+tmp[3542]*kernel[7]+tmp[3543]*kernel[8];
				ans[3443]<=tmp[3342]*kernel[0]+tmp[3343]*kernel[1]+tmp[3344]*kernel[2]+tmp[3442]*kernel[3]+tmp[3443]*kernel[4]+tmp[3444]*kernel[5]+tmp[3542]*kernel[6]+tmp[3543]*kernel[7]+tmp[3544]*kernel[8];
				ans[3444]<=tmp[3343]*kernel[0]+tmp[3344]*kernel[1]+tmp[3345]*kernel[2]+tmp[3443]*kernel[3]+tmp[3444]*kernel[4]+tmp[3445]*kernel[5]+tmp[3543]*kernel[6]+tmp[3544]*kernel[7]+tmp[3545]*kernel[8];
				ans[3445]<=tmp[3344]*kernel[0]+tmp[3345]*kernel[1]+tmp[3346]*kernel[2]+tmp[3444]*kernel[3]+tmp[3445]*kernel[4]+tmp[3446]*kernel[5]+tmp[3544]*kernel[6]+tmp[3545]*kernel[7]+tmp[3546]*kernel[8];
				ans[3446]<=tmp[3345]*kernel[0]+tmp[3346]*kernel[1]+tmp[3347]*kernel[2]+tmp[3445]*kernel[3]+tmp[3446]*kernel[4]+tmp[3447]*kernel[5]+tmp[3545]*kernel[6]+tmp[3546]*kernel[7]+tmp[3547]*kernel[8];
				ans[3447]<=tmp[3346]*kernel[0]+tmp[3347]*kernel[1]+tmp[3348]*kernel[2]+tmp[3446]*kernel[3]+tmp[3447]*kernel[4]+tmp[3448]*kernel[5]+tmp[3546]*kernel[6]+tmp[3547]*kernel[7]+tmp[3548]*kernel[8];
				ans[3448]<=tmp[3347]*kernel[0]+tmp[3348]*kernel[1]+tmp[3349]*kernel[2]+tmp[3447]*kernel[3]+tmp[3448]*kernel[4]+tmp[3449]*kernel[5]+tmp[3547]*kernel[6]+tmp[3548]*kernel[7]+tmp[3549]*kernel[8];
				ans[3449]<=tmp[3348]*kernel[0]+tmp[3349]*kernel[1]+tmp[3350]*kernel[2]+tmp[3448]*kernel[3]+tmp[3449]*kernel[4]+tmp[3450]*kernel[5]+tmp[3548]*kernel[6]+tmp[3549]*kernel[7]+tmp[3550]*kernel[8];
				ans[3450]<=tmp[3349]*kernel[0]+tmp[3350]*kernel[1]+tmp[3351]*kernel[2]+tmp[3449]*kernel[3]+tmp[3450]*kernel[4]+tmp[3451]*kernel[5]+tmp[3549]*kernel[6]+tmp[3550]*kernel[7]+tmp[3551]*kernel[8];
				ans[3451]<=tmp[3350]*kernel[0]+tmp[3351]*kernel[1]+tmp[3352]*kernel[2]+tmp[3450]*kernel[3]+tmp[3451]*kernel[4]+tmp[3452]*kernel[5]+tmp[3550]*kernel[6]+tmp[3551]*kernel[7]+tmp[3552]*kernel[8];
				ans[3452]<=tmp[3351]*kernel[0]+tmp[3352]*kernel[1]+tmp[3353]*kernel[2]+tmp[3451]*kernel[3]+tmp[3452]*kernel[4]+tmp[3453]*kernel[5]+tmp[3551]*kernel[6]+tmp[3552]*kernel[7]+tmp[3553]*kernel[8];
				ans[3453]<=tmp[3352]*kernel[0]+tmp[3353]*kernel[1]+tmp[3354]*kernel[2]+tmp[3452]*kernel[3]+tmp[3453]*kernel[4]+tmp[3454]*kernel[5]+tmp[3552]*kernel[6]+tmp[3553]*kernel[7]+tmp[3554]*kernel[8];
				ans[3454]<=tmp[3353]*kernel[0]+tmp[3354]*kernel[1]+tmp[3355]*kernel[2]+tmp[3453]*kernel[3]+tmp[3454]*kernel[4]+tmp[3455]*kernel[5]+tmp[3553]*kernel[6]+tmp[3554]*kernel[7]+tmp[3555]*kernel[8];
				ans[3455]<=tmp[3354]*kernel[0]+tmp[3355]*kernel[1]+tmp[3356]*kernel[2]+tmp[3454]*kernel[3]+tmp[3455]*kernel[4]+tmp[3456]*kernel[5]+tmp[3554]*kernel[6]+tmp[3555]*kernel[7]+tmp[3556]*kernel[8];
				ans[3456]<=tmp[3355]*kernel[0]+tmp[3356]*kernel[1]+tmp[3357]*kernel[2]+tmp[3455]*kernel[3]+tmp[3456]*kernel[4]+tmp[3457]*kernel[5]+tmp[3555]*kernel[6]+tmp[3556]*kernel[7]+tmp[3557]*kernel[8];
				ans[3457]<=tmp[3356]*kernel[0]+tmp[3357]*kernel[1]+tmp[3358]*kernel[2]+tmp[3456]*kernel[3]+tmp[3457]*kernel[4]+tmp[3458]*kernel[5]+tmp[3556]*kernel[6]+tmp[3557]*kernel[7]+tmp[3558]*kernel[8];
				ans[3458]<=tmp[3357]*kernel[0]+tmp[3358]*kernel[1]+tmp[3359]*kernel[2]+tmp[3457]*kernel[3]+tmp[3458]*kernel[4]+tmp[3459]*kernel[5]+tmp[3557]*kernel[6]+tmp[3558]*kernel[7]+tmp[3559]*kernel[8];
				ans[3459]<=tmp[3358]*kernel[0]+tmp[3359]*kernel[1]+tmp[3360]*kernel[2]+tmp[3458]*kernel[3]+tmp[3459]*kernel[4]+tmp[3460]*kernel[5]+tmp[3558]*kernel[6]+tmp[3559]*kernel[7]+tmp[3560]*kernel[8];
				ans[3460]<=tmp[3359]*kernel[0]+tmp[3360]*kernel[1]+tmp[3361]*kernel[2]+tmp[3459]*kernel[3]+tmp[3460]*kernel[4]+tmp[3461]*kernel[5]+tmp[3559]*kernel[6]+tmp[3560]*kernel[7]+tmp[3561]*kernel[8];
				ans[3461]<=tmp[3360]*kernel[0]+tmp[3361]*kernel[1]+tmp[3362]*kernel[2]+tmp[3460]*kernel[3]+tmp[3461]*kernel[4]+tmp[3462]*kernel[5]+tmp[3560]*kernel[6]+tmp[3561]*kernel[7]+tmp[3562]*kernel[8];
				ans[3462]<=tmp[3361]*kernel[0]+tmp[3362]*kernel[1]+tmp[3363]*kernel[2]+tmp[3461]*kernel[3]+tmp[3462]*kernel[4]+tmp[3463]*kernel[5]+tmp[3561]*kernel[6]+tmp[3562]*kernel[7]+tmp[3563]*kernel[8];
				ans[3463]<=tmp[3362]*kernel[0]+tmp[3363]*kernel[1]+tmp[3364]*kernel[2]+tmp[3462]*kernel[3]+tmp[3463]*kernel[4]+tmp[3464]*kernel[5]+tmp[3562]*kernel[6]+tmp[3563]*kernel[7]+tmp[3564]*kernel[8];
				ans[3464]<=tmp[3363]*kernel[0]+tmp[3364]*kernel[1]+tmp[3365]*kernel[2]+tmp[3463]*kernel[3]+tmp[3464]*kernel[4]+tmp[3465]*kernel[5]+tmp[3563]*kernel[6]+tmp[3564]*kernel[7]+tmp[3565]*kernel[8];
				ans[3465]<=tmp[3364]*kernel[0]+tmp[3365]*kernel[1]+tmp[3366]*kernel[2]+tmp[3464]*kernel[3]+tmp[3465]*kernel[4]+tmp[3466]*kernel[5]+tmp[3564]*kernel[6]+tmp[3565]*kernel[7]+tmp[3566]*kernel[8];
				ans[3466]<=tmp[3365]*kernel[0]+tmp[3366]*kernel[1]+tmp[3367]*kernel[2]+tmp[3465]*kernel[3]+tmp[3466]*kernel[4]+tmp[3467]*kernel[5]+tmp[3565]*kernel[6]+tmp[3566]*kernel[7]+tmp[3567]*kernel[8];
				ans[3467]<=tmp[3366]*kernel[0]+tmp[3367]*kernel[1]+tmp[3368]*kernel[2]+tmp[3466]*kernel[3]+tmp[3467]*kernel[4]+tmp[3468]*kernel[5]+tmp[3566]*kernel[6]+tmp[3567]*kernel[7]+tmp[3568]*kernel[8];
				ans[3468]<=tmp[3367]*kernel[0]+tmp[3368]*kernel[1]+tmp[3369]*kernel[2]+tmp[3467]*kernel[3]+tmp[3468]*kernel[4]+tmp[3469]*kernel[5]+tmp[3567]*kernel[6]+tmp[3568]*kernel[7]+tmp[3569]*kernel[8];
				ans[3469]<=tmp[3368]*kernel[0]+tmp[3369]*kernel[1]+tmp[3370]*kernel[2]+tmp[3468]*kernel[3]+tmp[3469]*kernel[4]+tmp[3470]*kernel[5]+tmp[3568]*kernel[6]+tmp[3569]*kernel[7]+tmp[3570]*kernel[8];
				ans[3470]<=tmp[3369]*kernel[0]+tmp[3370]*kernel[1]+tmp[3371]*kernel[2]+tmp[3469]*kernel[3]+tmp[3470]*kernel[4]+tmp[3471]*kernel[5]+tmp[3569]*kernel[6]+tmp[3570]*kernel[7]+tmp[3571]*kernel[8];
				ans[3471]<=tmp[3370]*kernel[0]+tmp[3371]*kernel[1]+tmp[3372]*kernel[2]+tmp[3470]*kernel[3]+tmp[3471]*kernel[4]+tmp[3472]*kernel[5]+tmp[3570]*kernel[6]+tmp[3571]*kernel[7]+tmp[3572]*kernel[8];
				ans[3472]<=tmp[3371]*kernel[0]+tmp[3372]*kernel[1]+tmp[3373]*kernel[2]+tmp[3471]*kernel[3]+tmp[3472]*kernel[4]+tmp[3473]*kernel[5]+tmp[3571]*kernel[6]+tmp[3572]*kernel[7]+tmp[3573]*kernel[8];
				ans[3473]<=tmp[3372]*kernel[0]+tmp[3373]*kernel[1]+tmp[3374]*kernel[2]+tmp[3472]*kernel[3]+tmp[3473]*kernel[4]+tmp[3474]*kernel[5]+tmp[3572]*kernel[6]+tmp[3573]*kernel[7]+tmp[3574]*kernel[8];
				ans[3474]<=tmp[3373]*kernel[0]+tmp[3374]*kernel[1]+tmp[3375]*kernel[2]+tmp[3473]*kernel[3]+tmp[3474]*kernel[4]+tmp[3475]*kernel[5]+tmp[3573]*kernel[6]+tmp[3574]*kernel[7]+tmp[3575]*kernel[8];
				ans[3475]<=tmp[3374]*kernel[0]+tmp[3375]*kernel[1]+tmp[3376]*kernel[2]+tmp[3474]*kernel[3]+tmp[3475]*kernel[4]+tmp[3476]*kernel[5]+tmp[3574]*kernel[6]+tmp[3575]*kernel[7]+tmp[3576]*kernel[8];
				ans[3476]<=tmp[3375]*kernel[0]+tmp[3376]*kernel[1]+tmp[3377]*kernel[2]+tmp[3475]*kernel[3]+tmp[3476]*kernel[4]+tmp[3477]*kernel[5]+tmp[3575]*kernel[6]+tmp[3576]*kernel[7]+tmp[3577]*kernel[8];
				ans[3477]<=tmp[3376]*kernel[0]+tmp[3377]*kernel[1]+tmp[3378]*kernel[2]+tmp[3476]*kernel[3]+tmp[3477]*kernel[4]+tmp[3478]*kernel[5]+tmp[3576]*kernel[6]+tmp[3577]*kernel[7]+tmp[3578]*kernel[8];
				ans[3478]<=tmp[3377]*kernel[0]+tmp[3378]*kernel[1]+tmp[3379]*kernel[2]+tmp[3477]*kernel[3]+tmp[3478]*kernel[4]+tmp[3479]*kernel[5]+tmp[3577]*kernel[6]+tmp[3578]*kernel[7]+tmp[3579]*kernel[8];
				ans[3479]<=tmp[3378]*kernel[0]+tmp[3379]*kernel[1]+tmp[3380]*kernel[2]+tmp[3478]*kernel[3]+tmp[3479]*kernel[4]+tmp[3480]*kernel[5]+tmp[3578]*kernel[6]+tmp[3579]*kernel[7]+tmp[3580]*kernel[8];
				ans[3480]<=tmp[3379]*kernel[0]+tmp[3380]*kernel[1]+tmp[3381]*kernel[2]+tmp[3479]*kernel[3]+tmp[3480]*kernel[4]+tmp[3481]*kernel[5]+tmp[3579]*kernel[6]+tmp[3580]*kernel[7]+tmp[3581]*kernel[8];
				ans[3481]<=tmp[3380]*kernel[0]+tmp[3381]*kernel[1]+tmp[3382]*kernel[2]+tmp[3480]*kernel[3]+tmp[3481]*kernel[4]+tmp[3482]*kernel[5]+tmp[3580]*kernel[6]+tmp[3581]*kernel[7]+tmp[3582]*kernel[8];
				ans[3482]<=tmp[3381]*kernel[0]+tmp[3382]*kernel[1]+tmp[3383]*kernel[2]+tmp[3481]*kernel[3]+tmp[3482]*kernel[4]+tmp[3483]*kernel[5]+tmp[3581]*kernel[6]+tmp[3582]*kernel[7]+tmp[3583]*kernel[8];
				ans[3483]<=tmp[3382]*kernel[0]+tmp[3383]*kernel[1]+tmp[3384]*kernel[2]+tmp[3482]*kernel[3]+tmp[3483]*kernel[4]+tmp[3484]*kernel[5]+tmp[3582]*kernel[6]+tmp[3583]*kernel[7]+tmp[3584]*kernel[8];
				ans[3484]<=tmp[3383]*kernel[0]+tmp[3384]*kernel[1]+tmp[3385]*kernel[2]+tmp[3483]*kernel[3]+tmp[3484]*kernel[4]+tmp[3485]*kernel[5]+tmp[3583]*kernel[6]+tmp[3584]*kernel[7]+tmp[3585]*kernel[8];
				ans[3485]<=tmp[3384]*kernel[0]+tmp[3385]*kernel[1]+tmp[3386]*kernel[2]+tmp[3484]*kernel[3]+tmp[3485]*kernel[4]+tmp[3486]*kernel[5]+tmp[3584]*kernel[6]+tmp[3585]*kernel[7]+tmp[3586]*kernel[8];
				ans[3486]<=tmp[3385]*kernel[0]+tmp[3386]*kernel[1]+tmp[3387]*kernel[2]+tmp[3485]*kernel[3]+tmp[3486]*kernel[4]+tmp[3487]*kernel[5]+tmp[3585]*kernel[6]+tmp[3586]*kernel[7]+tmp[3587]*kernel[8];
				ans[3487]<=tmp[3386]*kernel[0]+tmp[3387]*kernel[1]+tmp[3388]*kernel[2]+tmp[3486]*kernel[3]+tmp[3487]*kernel[4]+tmp[3488]*kernel[5]+tmp[3586]*kernel[6]+tmp[3587]*kernel[7]+tmp[3588]*kernel[8];
				ans[3488]<=tmp[3387]*kernel[0]+tmp[3388]*kernel[1]+tmp[3389]*kernel[2]+tmp[3487]*kernel[3]+tmp[3488]*kernel[4]+tmp[3489]*kernel[5]+tmp[3587]*kernel[6]+tmp[3588]*kernel[7]+tmp[3589]*kernel[8];
				ans[3489]<=tmp[3388]*kernel[0]+tmp[3389]*kernel[1]+tmp[3390]*kernel[2]+tmp[3488]*kernel[3]+tmp[3489]*kernel[4]+tmp[3490]*kernel[5]+tmp[3588]*kernel[6]+tmp[3589]*kernel[7]+tmp[3590]*kernel[8];
				ans[3490]<=tmp[3389]*kernel[0]+tmp[3390]*kernel[1]+tmp[3391]*kernel[2]+tmp[3489]*kernel[3]+tmp[3490]*kernel[4]+tmp[3491]*kernel[5]+tmp[3589]*kernel[6]+tmp[3590]*kernel[7]+tmp[3591]*kernel[8];
				ans[3491]<=tmp[3390]*kernel[0]+tmp[3391]*kernel[1]+tmp[3392]*kernel[2]+tmp[3490]*kernel[3]+tmp[3491]*kernel[4]+tmp[3492]*kernel[5]+tmp[3590]*kernel[6]+tmp[3591]*kernel[7]+tmp[3592]*kernel[8];
				ans[3492]<=tmp[3391]*kernel[0]+tmp[3392]*kernel[1]+tmp[3393]*kernel[2]+tmp[3491]*kernel[3]+tmp[3492]*kernel[4]+tmp[3493]*kernel[5]+tmp[3591]*kernel[6]+tmp[3592]*kernel[7]+tmp[3593]*kernel[8];
				ans[3493]<=tmp[3392]*kernel[0]+tmp[3393]*kernel[1]+tmp[3394]*kernel[2]+tmp[3492]*kernel[3]+tmp[3493]*kernel[4]+tmp[3494]*kernel[5]+tmp[3592]*kernel[6]+tmp[3593]*kernel[7]+tmp[3594]*kernel[8];
				ans[3494]<=tmp[3393]*kernel[0]+tmp[3394]*kernel[1]+tmp[3395]*kernel[2]+tmp[3493]*kernel[3]+tmp[3494]*kernel[4]+tmp[3495]*kernel[5]+tmp[3593]*kernel[6]+tmp[3594]*kernel[7]+tmp[3595]*kernel[8];
				ans[3495]<=tmp[3394]*kernel[0]+tmp[3395]*kernel[1]+tmp[3396]*kernel[2]+tmp[3494]*kernel[3]+tmp[3495]*kernel[4]+tmp[3496]*kernel[5]+tmp[3594]*kernel[6]+tmp[3595]*kernel[7]+tmp[3596]*kernel[8];
				ans[3496]<=tmp[3395]*kernel[0]+tmp[3396]*kernel[1]+tmp[3397]*kernel[2]+tmp[3495]*kernel[3]+tmp[3496]*kernel[4]+tmp[3497]*kernel[5]+tmp[3595]*kernel[6]+tmp[3596]*kernel[7]+tmp[3597]*kernel[8];
				ans[3497]<=tmp[3396]*kernel[0]+tmp[3397]*kernel[1]+tmp[3398]*kernel[2]+tmp[3496]*kernel[3]+tmp[3497]*kernel[4]+tmp[3498]*kernel[5]+tmp[3596]*kernel[6]+tmp[3597]*kernel[7]+tmp[3598]*kernel[8];
				ans[3498]<=tmp[3397]*kernel[0]+tmp[3398]*kernel[1]+tmp[3399]*kernel[2]+tmp[3497]*kernel[3]+tmp[3498]*kernel[4]+tmp[3499]*kernel[5]+tmp[3597]*kernel[6]+tmp[3598]*kernel[7]+tmp[3599]*kernel[8];
				ans[3499]<=tmp[3398]*kernel[0]+tmp[3399]*kernel[1]+tmp[3498]*kernel[3]+tmp[3499]*kernel[4]+tmp[3598]*kernel[6]+tmp[3599]*kernel[7];
				ans[3500]<=tmp[3400]*kernel[1]+tmp[3401]*kernel[2]+tmp[3500]*kernel[4]+tmp[3501]*kernel[5]+tmp[3600]*kernel[7]+tmp[3601]*kernel[8];
				ans[3501]<=tmp[3400]*kernel[0]+tmp[3401]*kernel[1]+tmp[3402]*kernel[2]+tmp[3500]*kernel[3]+tmp[3501]*kernel[4]+tmp[3502]*kernel[5]+tmp[3600]*kernel[6]+tmp[3601]*kernel[7]+tmp[3602]*kernel[8];
				ans[3502]<=tmp[3401]*kernel[0]+tmp[3402]*kernel[1]+tmp[3403]*kernel[2]+tmp[3501]*kernel[3]+tmp[3502]*kernel[4]+tmp[3503]*kernel[5]+tmp[3601]*kernel[6]+tmp[3602]*kernel[7]+tmp[3603]*kernel[8];
				ans[3503]<=tmp[3402]*kernel[0]+tmp[3403]*kernel[1]+tmp[3404]*kernel[2]+tmp[3502]*kernel[3]+tmp[3503]*kernel[4]+tmp[3504]*kernel[5]+tmp[3602]*kernel[6]+tmp[3603]*kernel[7]+tmp[3604]*kernel[8];
				ans[3504]<=tmp[3403]*kernel[0]+tmp[3404]*kernel[1]+tmp[3405]*kernel[2]+tmp[3503]*kernel[3]+tmp[3504]*kernel[4]+tmp[3505]*kernel[5]+tmp[3603]*kernel[6]+tmp[3604]*kernel[7]+tmp[3605]*kernel[8];
				ans[3505]<=tmp[3404]*kernel[0]+tmp[3405]*kernel[1]+tmp[3406]*kernel[2]+tmp[3504]*kernel[3]+tmp[3505]*kernel[4]+tmp[3506]*kernel[5]+tmp[3604]*kernel[6]+tmp[3605]*kernel[7]+tmp[3606]*kernel[8];
				ans[3506]<=tmp[3405]*kernel[0]+tmp[3406]*kernel[1]+tmp[3407]*kernel[2]+tmp[3505]*kernel[3]+tmp[3506]*kernel[4]+tmp[3507]*kernel[5]+tmp[3605]*kernel[6]+tmp[3606]*kernel[7]+tmp[3607]*kernel[8];
				ans[3507]<=tmp[3406]*kernel[0]+tmp[3407]*kernel[1]+tmp[3408]*kernel[2]+tmp[3506]*kernel[3]+tmp[3507]*kernel[4]+tmp[3508]*kernel[5]+tmp[3606]*kernel[6]+tmp[3607]*kernel[7]+tmp[3608]*kernel[8];
				ans[3508]<=tmp[3407]*kernel[0]+tmp[3408]*kernel[1]+tmp[3409]*kernel[2]+tmp[3507]*kernel[3]+tmp[3508]*kernel[4]+tmp[3509]*kernel[5]+tmp[3607]*kernel[6]+tmp[3608]*kernel[7]+tmp[3609]*kernel[8];
				ans[3509]<=tmp[3408]*kernel[0]+tmp[3409]*kernel[1]+tmp[3410]*kernel[2]+tmp[3508]*kernel[3]+tmp[3509]*kernel[4]+tmp[3510]*kernel[5]+tmp[3608]*kernel[6]+tmp[3609]*kernel[7]+tmp[3610]*kernel[8];
				ans[3510]<=tmp[3409]*kernel[0]+tmp[3410]*kernel[1]+tmp[3411]*kernel[2]+tmp[3509]*kernel[3]+tmp[3510]*kernel[4]+tmp[3511]*kernel[5]+tmp[3609]*kernel[6]+tmp[3610]*kernel[7]+tmp[3611]*kernel[8];
				ans[3511]<=tmp[3410]*kernel[0]+tmp[3411]*kernel[1]+tmp[3412]*kernel[2]+tmp[3510]*kernel[3]+tmp[3511]*kernel[4]+tmp[3512]*kernel[5]+tmp[3610]*kernel[6]+tmp[3611]*kernel[7]+tmp[3612]*kernel[8];
				ans[3512]<=tmp[3411]*kernel[0]+tmp[3412]*kernel[1]+tmp[3413]*kernel[2]+tmp[3511]*kernel[3]+tmp[3512]*kernel[4]+tmp[3513]*kernel[5]+tmp[3611]*kernel[6]+tmp[3612]*kernel[7]+tmp[3613]*kernel[8];
				ans[3513]<=tmp[3412]*kernel[0]+tmp[3413]*kernel[1]+tmp[3414]*kernel[2]+tmp[3512]*kernel[3]+tmp[3513]*kernel[4]+tmp[3514]*kernel[5]+tmp[3612]*kernel[6]+tmp[3613]*kernel[7]+tmp[3614]*kernel[8];
				ans[3514]<=tmp[3413]*kernel[0]+tmp[3414]*kernel[1]+tmp[3415]*kernel[2]+tmp[3513]*kernel[3]+tmp[3514]*kernel[4]+tmp[3515]*kernel[5]+tmp[3613]*kernel[6]+tmp[3614]*kernel[7]+tmp[3615]*kernel[8];
				ans[3515]<=tmp[3414]*kernel[0]+tmp[3415]*kernel[1]+tmp[3416]*kernel[2]+tmp[3514]*kernel[3]+tmp[3515]*kernel[4]+tmp[3516]*kernel[5]+tmp[3614]*kernel[6]+tmp[3615]*kernel[7]+tmp[3616]*kernel[8];
				ans[3516]<=tmp[3415]*kernel[0]+tmp[3416]*kernel[1]+tmp[3417]*kernel[2]+tmp[3515]*kernel[3]+tmp[3516]*kernel[4]+tmp[3517]*kernel[5]+tmp[3615]*kernel[6]+tmp[3616]*kernel[7]+tmp[3617]*kernel[8];
				ans[3517]<=tmp[3416]*kernel[0]+tmp[3417]*kernel[1]+tmp[3418]*kernel[2]+tmp[3516]*kernel[3]+tmp[3517]*kernel[4]+tmp[3518]*kernel[5]+tmp[3616]*kernel[6]+tmp[3617]*kernel[7]+tmp[3618]*kernel[8];
				ans[3518]<=tmp[3417]*kernel[0]+tmp[3418]*kernel[1]+tmp[3419]*kernel[2]+tmp[3517]*kernel[3]+tmp[3518]*kernel[4]+tmp[3519]*kernel[5]+tmp[3617]*kernel[6]+tmp[3618]*kernel[7]+tmp[3619]*kernel[8];
				ans[3519]<=tmp[3418]*kernel[0]+tmp[3419]*kernel[1]+tmp[3420]*kernel[2]+tmp[3518]*kernel[3]+tmp[3519]*kernel[4]+tmp[3520]*kernel[5]+tmp[3618]*kernel[6]+tmp[3619]*kernel[7]+tmp[3620]*kernel[8];
				ans[3520]<=tmp[3419]*kernel[0]+tmp[3420]*kernel[1]+tmp[3421]*kernel[2]+tmp[3519]*kernel[3]+tmp[3520]*kernel[4]+tmp[3521]*kernel[5]+tmp[3619]*kernel[6]+tmp[3620]*kernel[7]+tmp[3621]*kernel[8];
				ans[3521]<=tmp[3420]*kernel[0]+tmp[3421]*kernel[1]+tmp[3422]*kernel[2]+tmp[3520]*kernel[3]+tmp[3521]*kernel[4]+tmp[3522]*kernel[5]+tmp[3620]*kernel[6]+tmp[3621]*kernel[7]+tmp[3622]*kernel[8];
				ans[3522]<=tmp[3421]*kernel[0]+tmp[3422]*kernel[1]+tmp[3423]*kernel[2]+tmp[3521]*kernel[3]+tmp[3522]*kernel[4]+tmp[3523]*kernel[5]+tmp[3621]*kernel[6]+tmp[3622]*kernel[7]+tmp[3623]*kernel[8];
				ans[3523]<=tmp[3422]*kernel[0]+tmp[3423]*kernel[1]+tmp[3424]*kernel[2]+tmp[3522]*kernel[3]+tmp[3523]*kernel[4]+tmp[3524]*kernel[5]+tmp[3622]*kernel[6]+tmp[3623]*kernel[7]+tmp[3624]*kernel[8];
				ans[3524]<=tmp[3423]*kernel[0]+tmp[3424]*kernel[1]+tmp[3425]*kernel[2]+tmp[3523]*kernel[3]+tmp[3524]*kernel[4]+tmp[3525]*kernel[5]+tmp[3623]*kernel[6]+tmp[3624]*kernel[7]+tmp[3625]*kernel[8];
				ans[3525]<=tmp[3424]*kernel[0]+tmp[3425]*kernel[1]+tmp[3426]*kernel[2]+tmp[3524]*kernel[3]+tmp[3525]*kernel[4]+tmp[3526]*kernel[5]+tmp[3624]*kernel[6]+tmp[3625]*kernel[7]+tmp[3626]*kernel[8];
				ans[3526]<=tmp[3425]*kernel[0]+tmp[3426]*kernel[1]+tmp[3427]*kernel[2]+tmp[3525]*kernel[3]+tmp[3526]*kernel[4]+tmp[3527]*kernel[5]+tmp[3625]*kernel[6]+tmp[3626]*kernel[7]+tmp[3627]*kernel[8];
				ans[3527]<=tmp[3426]*kernel[0]+tmp[3427]*kernel[1]+tmp[3428]*kernel[2]+tmp[3526]*kernel[3]+tmp[3527]*kernel[4]+tmp[3528]*kernel[5]+tmp[3626]*kernel[6]+tmp[3627]*kernel[7]+tmp[3628]*kernel[8];
				ans[3528]<=tmp[3427]*kernel[0]+tmp[3428]*kernel[1]+tmp[3429]*kernel[2]+tmp[3527]*kernel[3]+tmp[3528]*kernel[4]+tmp[3529]*kernel[5]+tmp[3627]*kernel[6]+tmp[3628]*kernel[7]+tmp[3629]*kernel[8];
				ans[3529]<=tmp[3428]*kernel[0]+tmp[3429]*kernel[1]+tmp[3430]*kernel[2]+tmp[3528]*kernel[3]+tmp[3529]*kernel[4]+tmp[3530]*kernel[5]+tmp[3628]*kernel[6]+tmp[3629]*kernel[7]+tmp[3630]*kernel[8];
				ans[3530]<=tmp[3429]*kernel[0]+tmp[3430]*kernel[1]+tmp[3431]*kernel[2]+tmp[3529]*kernel[3]+tmp[3530]*kernel[4]+tmp[3531]*kernel[5]+tmp[3629]*kernel[6]+tmp[3630]*kernel[7]+tmp[3631]*kernel[8];
				ans[3531]<=tmp[3430]*kernel[0]+tmp[3431]*kernel[1]+tmp[3432]*kernel[2]+tmp[3530]*kernel[3]+tmp[3531]*kernel[4]+tmp[3532]*kernel[5]+tmp[3630]*kernel[6]+tmp[3631]*kernel[7]+tmp[3632]*kernel[8];
				ans[3532]<=tmp[3431]*kernel[0]+tmp[3432]*kernel[1]+tmp[3433]*kernel[2]+tmp[3531]*kernel[3]+tmp[3532]*kernel[4]+tmp[3533]*kernel[5]+tmp[3631]*kernel[6]+tmp[3632]*kernel[7]+tmp[3633]*kernel[8];
				ans[3533]<=tmp[3432]*kernel[0]+tmp[3433]*kernel[1]+tmp[3434]*kernel[2]+tmp[3532]*kernel[3]+tmp[3533]*kernel[4]+tmp[3534]*kernel[5]+tmp[3632]*kernel[6]+tmp[3633]*kernel[7]+tmp[3634]*kernel[8];
				ans[3534]<=tmp[3433]*kernel[0]+tmp[3434]*kernel[1]+tmp[3435]*kernel[2]+tmp[3533]*kernel[3]+tmp[3534]*kernel[4]+tmp[3535]*kernel[5]+tmp[3633]*kernel[6]+tmp[3634]*kernel[7]+tmp[3635]*kernel[8];
				ans[3535]<=tmp[3434]*kernel[0]+tmp[3435]*kernel[1]+tmp[3436]*kernel[2]+tmp[3534]*kernel[3]+tmp[3535]*kernel[4]+tmp[3536]*kernel[5]+tmp[3634]*kernel[6]+tmp[3635]*kernel[7]+tmp[3636]*kernel[8];
				ans[3536]<=tmp[3435]*kernel[0]+tmp[3436]*kernel[1]+tmp[3437]*kernel[2]+tmp[3535]*kernel[3]+tmp[3536]*kernel[4]+tmp[3537]*kernel[5]+tmp[3635]*kernel[6]+tmp[3636]*kernel[7]+tmp[3637]*kernel[8];
				ans[3537]<=tmp[3436]*kernel[0]+tmp[3437]*kernel[1]+tmp[3438]*kernel[2]+tmp[3536]*kernel[3]+tmp[3537]*kernel[4]+tmp[3538]*kernel[5]+tmp[3636]*kernel[6]+tmp[3637]*kernel[7]+tmp[3638]*kernel[8];
				ans[3538]<=tmp[3437]*kernel[0]+tmp[3438]*kernel[1]+tmp[3439]*kernel[2]+tmp[3537]*kernel[3]+tmp[3538]*kernel[4]+tmp[3539]*kernel[5]+tmp[3637]*kernel[6]+tmp[3638]*kernel[7]+tmp[3639]*kernel[8];
				ans[3539]<=tmp[3438]*kernel[0]+tmp[3439]*kernel[1]+tmp[3440]*kernel[2]+tmp[3538]*kernel[3]+tmp[3539]*kernel[4]+tmp[3540]*kernel[5]+tmp[3638]*kernel[6]+tmp[3639]*kernel[7]+tmp[3640]*kernel[8];
				ans[3540]<=tmp[3439]*kernel[0]+tmp[3440]*kernel[1]+tmp[3441]*kernel[2]+tmp[3539]*kernel[3]+tmp[3540]*kernel[4]+tmp[3541]*kernel[5]+tmp[3639]*kernel[6]+tmp[3640]*kernel[7]+tmp[3641]*kernel[8];
				ans[3541]<=tmp[3440]*kernel[0]+tmp[3441]*kernel[1]+tmp[3442]*kernel[2]+tmp[3540]*kernel[3]+tmp[3541]*kernel[4]+tmp[3542]*kernel[5]+tmp[3640]*kernel[6]+tmp[3641]*kernel[7]+tmp[3642]*kernel[8];
				ans[3542]<=tmp[3441]*kernel[0]+tmp[3442]*kernel[1]+tmp[3443]*kernel[2]+tmp[3541]*kernel[3]+tmp[3542]*kernel[4]+tmp[3543]*kernel[5]+tmp[3641]*kernel[6]+tmp[3642]*kernel[7]+tmp[3643]*kernel[8];
				ans[3543]<=tmp[3442]*kernel[0]+tmp[3443]*kernel[1]+tmp[3444]*kernel[2]+tmp[3542]*kernel[3]+tmp[3543]*kernel[4]+tmp[3544]*kernel[5]+tmp[3642]*kernel[6]+tmp[3643]*kernel[7]+tmp[3644]*kernel[8];
				ans[3544]<=tmp[3443]*kernel[0]+tmp[3444]*kernel[1]+tmp[3445]*kernel[2]+tmp[3543]*kernel[3]+tmp[3544]*kernel[4]+tmp[3545]*kernel[5]+tmp[3643]*kernel[6]+tmp[3644]*kernel[7]+tmp[3645]*kernel[8];
				ans[3545]<=tmp[3444]*kernel[0]+tmp[3445]*kernel[1]+tmp[3446]*kernel[2]+tmp[3544]*kernel[3]+tmp[3545]*kernel[4]+tmp[3546]*kernel[5]+tmp[3644]*kernel[6]+tmp[3645]*kernel[7]+tmp[3646]*kernel[8];
				ans[3546]<=tmp[3445]*kernel[0]+tmp[3446]*kernel[1]+tmp[3447]*kernel[2]+tmp[3545]*kernel[3]+tmp[3546]*kernel[4]+tmp[3547]*kernel[5]+tmp[3645]*kernel[6]+tmp[3646]*kernel[7]+tmp[3647]*kernel[8];
				ans[3547]<=tmp[3446]*kernel[0]+tmp[3447]*kernel[1]+tmp[3448]*kernel[2]+tmp[3546]*kernel[3]+tmp[3547]*kernel[4]+tmp[3548]*kernel[5]+tmp[3646]*kernel[6]+tmp[3647]*kernel[7]+tmp[3648]*kernel[8];
				ans[3548]<=tmp[3447]*kernel[0]+tmp[3448]*kernel[1]+tmp[3449]*kernel[2]+tmp[3547]*kernel[3]+tmp[3548]*kernel[4]+tmp[3549]*kernel[5]+tmp[3647]*kernel[6]+tmp[3648]*kernel[7]+tmp[3649]*kernel[8];
				ans[3549]<=tmp[3448]*kernel[0]+tmp[3449]*kernel[1]+tmp[3450]*kernel[2]+tmp[3548]*kernel[3]+tmp[3549]*kernel[4]+tmp[3550]*kernel[5]+tmp[3648]*kernel[6]+tmp[3649]*kernel[7]+tmp[3650]*kernel[8];
				ans[3550]<=tmp[3449]*kernel[0]+tmp[3450]*kernel[1]+tmp[3451]*kernel[2]+tmp[3549]*kernel[3]+tmp[3550]*kernel[4]+tmp[3551]*kernel[5]+tmp[3649]*kernel[6]+tmp[3650]*kernel[7]+tmp[3651]*kernel[8];
				ans[3551]<=tmp[3450]*kernel[0]+tmp[3451]*kernel[1]+tmp[3452]*kernel[2]+tmp[3550]*kernel[3]+tmp[3551]*kernel[4]+tmp[3552]*kernel[5]+tmp[3650]*kernel[6]+tmp[3651]*kernel[7]+tmp[3652]*kernel[8];
				ans[3552]<=tmp[3451]*kernel[0]+tmp[3452]*kernel[1]+tmp[3453]*kernel[2]+tmp[3551]*kernel[3]+tmp[3552]*kernel[4]+tmp[3553]*kernel[5]+tmp[3651]*kernel[6]+tmp[3652]*kernel[7]+tmp[3653]*kernel[8];
				ans[3553]<=tmp[3452]*kernel[0]+tmp[3453]*kernel[1]+tmp[3454]*kernel[2]+tmp[3552]*kernel[3]+tmp[3553]*kernel[4]+tmp[3554]*kernel[5]+tmp[3652]*kernel[6]+tmp[3653]*kernel[7]+tmp[3654]*kernel[8];
				ans[3554]<=tmp[3453]*kernel[0]+tmp[3454]*kernel[1]+tmp[3455]*kernel[2]+tmp[3553]*kernel[3]+tmp[3554]*kernel[4]+tmp[3555]*kernel[5]+tmp[3653]*kernel[6]+tmp[3654]*kernel[7]+tmp[3655]*kernel[8];
				ans[3555]<=tmp[3454]*kernel[0]+tmp[3455]*kernel[1]+tmp[3456]*kernel[2]+tmp[3554]*kernel[3]+tmp[3555]*kernel[4]+tmp[3556]*kernel[5]+tmp[3654]*kernel[6]+tmp[3655]*kernel[7]+tmp[3656]*kernel[8];
				ans[3556]<=tmp[3455]*kernel[0]+tmp[3456]*kernel[1]+tmp[3457]*kernel[2]+tmp[3555]*kernel[3]+tmp[3556]*kernel[4]+tmp[3557]*kernel[5]+tmp[3655]*kernel[6]+tmp[3656]*kernel[7]+tmp[3657]*kernel[8];
				ans[3557]<=tmp[3456]*kernel[0]+tmp[3457]*kernel[1]+tmp[3458]*kernel[2]+tmp[3556]*kernel[3]+tmp[3557]*kernel[4]+tmp[3558]*kernel[5]+tmp[3656]*kernel[6]+tmp[3657]*kernel[7]+tmp[3658]*kernel[8];
				ans[3558]<=tmp[3457]*kernel[0]+tmp[3458]*kernel[1]+tmp[3459]*kernel[2]+tmp[3557]*kernel[3]+tmp[3558]*kernel[4]+tmp[3559]*kernel[5]+tmp[3657]*kernel[6]+tmp[3658]*kernel[7]+tmp[3659]*kernel[8];
				ans[3559]<=tmp[3458]*kernel[0]+tmp[3459]*kernel[1]+tmp[3460]*kernel[2]+tmp[3558]*kernel[3]+tmp[3559]*kernel[4]+tmp[3560]*kernel[5]+tmp[3658]*kernel[6]+tmp[3659]*kernel[7]+tmp[3660]*kernel[8];
				ans[3560]<=tmp[3459]*kernel[0]+tmp[3460]*kernel[1]+tmp[3461]*kernel[2]+tmp[3559]*kernel[3]+tmp[3560]*kernel[4]+tmp[3561]*kernel[5]+tmp[3659]*kernel[6]+tmp[3660]*kernel[7]+tmp[3661]*kernel[8];
				ans[3561]<=tmp[3460]*kernel[0]+tmp[3461]*kernel[1]+tmp[3462]*kernel[2]+tmp[3560]*kernel[3]+tmp[3561]*kernel[4]+tmp[3562]*kernel[5]+tmp[3660]*kernel[6]+tmp[3661]*kernel[7]+tmp[3662]*kernel[8];
				ans[3562]<=tmp[3461]*kernel[0]+tmp[3462]*kernel[1]+tmp[3463]*kernel[2]+tmp[3561]*kernel[3]+tmp[3562]*kernel[4]+tmp[3563]*kernel[5]+tmp[3661]*kernel[6]+tmp[3662]*kernel[7]+tmp[3663]*kernel[8];
				ans[3563]<=tmp[3462]*kernel[0]+tmp[3463]*kernel[1]+tmp[3464]*kernel[2]+tmp[3562]*kernel[3]+tmp[3563]*kernel[4]+tmp[3564]*kernel[5]+tmp[3662]*kernel[6]+tmp[3663]*kernel[7]+tmp[3664]*kernel[8];
				ans[3564]<=tmp[3463]*kernel[0]+tmp[3464]*kernel[1]+tmp[3465]*kernel[2]+tmp[3563]*kernel[3]+tmp[3564]*kernel[4]+tmp[3565]*kernel[5]+tmp[3663]*kernel[6]+tmp[3664]*kernel[7]+tmp[3665]*kernel[8];
				ans[3565]<=tmp[3464]*kernel[0]+tmp[3465]*kernel[1]+tmp[3466]*kernel[2]+tmp[3564]*kernel[3]+tmp[3565]*kernel[4]+tmp[3566]*kernel[5]+tmp[3664]*kernel[6]+tmp[3665]*kernel[7]+tmp[3666]*kernel[8];
				ans[3566]<=tmp[3465]*kernel[0]+tmp[3466]*kernel[1]+tmp[3467]*kernel[2]+tmp[3565]*kernel[3]+tmp[3566]*kernel[4]+tmp[3567]*kernel[5]+tmp[3665]*kernel[6]+tmp[3666]*kernel[7]+tmp[3667]*kernel[8];
				ans[3567]<=tmp[3466]*kernel[0]+tmp[3467]*kernel[1]+tmp[3468]*kernel[2]+tmp[3566]*kernel[3]+tmp[3567]*kernel[4]+tmp[3568]*kernel[5]+tmp[3666]*kernel[6]+tmp[3667]*kernel[7]+tmp[3668]*kernel[8];
				ans[3568]<=tmp[3467]*kernel[0]+tmp[3468]*kernel[1]+tmp[3469]*kernel[2]+tmp[3567]*kernel[3]+tmp[3568]*kernel[4]+tmp[3569]*kernel[5]+tmp[3667]*kernel[6]+tmp[3668]*kernel[7]+tmp[3669]*kernel[8];
				ans[3569]<=tmp[3468]*kernel[0]+tmp[3469]*kernel[1]+tmp[3470]*kernel[2]+tmp[3568]*kernel[3]+tmp[3569]*kernel[4]+tmp[3570]*kernel[5]+tmp[3668]*kernel[6]+tmp[3669]*kernel[7]+tmp[3670]*kernel[8];
				ans[3570]<=tmp[3469]*kernel[0]+tmp[3470]*kernel[1]+tmp[3471]*kernel[2]+tmp[3569]*kernel[3]+tmp[3570]*kernel[4]+tmp[3571]*kernel[5]+tmp[3669]*kernel[6]+tmp[3670]*kernel[7]+tmp[3671]*kernel[8];
				ans[3571]<=tmp[3470]*kernel[0]+tmp[3471]*kernel[1]+tmp[3472]*kernel[2]+tmp[3570]*kernel[3]+tmp[3571]*kernel[4]+tmp[3572]*kernel[5]+tmp[3670]*kernel[6]+tmp[3671]*kernel[7]+tmp[3672]*kernel[8];
				ans[3572]<=tmp[3471]*kernel[0]+tmp[3472]*kernel[1]+tmp[3473]*kernel[2]+tmp[3571]*kernel[3]+tmp[3572]*kernel[4]+tmp[3573]*kernel[5]+tmp[3671]*kernel[6]+tmp[3672]*kernel[7]+tmp[3673]*kernel[8];
				ans[3573]<=tmp[3472]*kernel[0]+tmp[3473]*kernel[1]+tmp[3474]*kernel[2]+tmp[3572]*kernel[3]+tmp[3573]*kernel[4]+tmp[3574]*kernel[5]+tmp[3672]*kernel[6]+tmp[3673]*kernel[7]+tmp[3674]*kernel[8];
				ans[3574]<=tmp[3473]*kernel[0]+tmp[3474]*kernel[1]+tmp[3475]*kernel[2]+tmp[3573]*kernel[3]+tmp[3574]*kernel[4]+tmp[3575]*kernel[5]+tmp[3673]*kernel[6]+tmp[3674]*kernel[7]+tmp[3675]*kernel[8];
				ans[3575]<=tmp[3474]*kernel[0]+tmp[3475]*kernel[1]+tmp[3476]*kernel[2]+tmp[3574]*kernel[3]+tmp[3575]*kernel[4]+tmp[3576]*kernel[5]+tmp[3674]*kernel[6]+tmp[3675]*kernel[7]+tmp[3676]*kernel[8];
				ans[3576]<=tmp[3475]*kernel[0]+tmp[3476]*kernel[1]+tmp[3477]*kernel[2]+tmp[3575]*kernel[3]+tmp[3576]*kernel[4]+tmp[3577]*kernel[5]+tmp[3675]*kernel[6]+tmp[3676]*kernel[7]+tmp[3677]*kernel[8];
				ans[3577]<=tmp[3476]*kernel[0]+tmp[3477]*kernel[1]+tmp[3478]*kernel[2]+tmp[3576]*kernel[3]+tmp[3577]*kernel[4]+tmp[3578]*kernel[5]+tmp[3676]*kernel[6]+tmp[3677]*kernel[7]+tmp[3678]*kernel[8];
				ans[3578]<=tmp[3477]*kernel[0]+tmp[3478]*kernel[1]+tmp[3479]*kernel[2]+tmp[3577]*kernel[3]+tmp[3578]*kernel[4]+tmp[3579]*kernel[5]+tmp[3677]*kernel[6]+tmp[3678]*kernel[7]+tmp[3679]*kernel[8];
				ans[3579]<=tmp[3478]*kernel[0]+tmp[3479]*kernel[1]+tmp[3480]*kernel[2]+tmp[3578]*kernel[3]+tmp[3579]*kernel[4]+tmp[3580]*kernel[5]+tmp[3678]*kernel[6]+tmp[3679]*kernel[7]+tmp[3680]*kernel[8];
				ans[3580]<=tmp[3479]*kernel[0]+tmp[3480]*kernel[1]+tmp[3481]*kernel[2]+tmp[3579]*kernel[3]+tmp[3580]*kernel[4]+tmp[3581]*kernel[5]+tmp[3679]*kernel[6]+tmp[3680]*kernel[7]+tmp[3681]*kernel[8];
				ans[3581]<=tmp[3480]*kernel[0]+tmp[3481]*kernel[1]+tmp[3482]*kernel[2]+tmp[3580]*kernel[3]+tmp[3581]*kernel[4]+tmp[3582]*kernel[5]+tmp[3680]*kernel[6]+tmp[3681]*kernel[7]+tmp[3682]*kernel[8];
				ans[3582]<=tmp[3481]*kernel[0]+tmp[3482]*kernel[1]+tmp[3483]*kernel[2]+tmp[3581]*kernel[3]+tmp[3582]*kernel[4]+tmp[3583]*kernel[5]+tmp[3681]*kernel[6]+tmp[3682]*kernel[7]+tmp[3683]*kernel[8];
				ans[3583]<=tmp[3482]*kernel[0]+tmp[3483]*kernel[1]+tmp[3484]*kernel[2]+tmp[3582]*kernel[3]+tmp[3583]*kernel[4]+tmp[3584]*kernel[5]+tmp[3682]*kernel[6]+tmp[3683]*kernel[7]+tmp[3684]*kernel[8];
				ans[3584]<=tmp[3483]*kernel[0]+tmp[3484]*kernel[1]+tmp[3485]*kernel[2]+tmp[3583]*kernel[3]+tmp[3584]*kernel[4]+tmp[3585]*kernel[5]+tmp[3683]*kernel[6]+tmp[3684]*kernel[7]+tmp[3685]*kernel[8];
				ans[3585]<=tmp[3484]*kernel[0]+tmp[3485]*kernel[1]+tmp[3486]*kernel[2]+tmp[3584]*kernel[3]+tmp[3585]*kernel[4]+tmp[3586]*kernel[5]+tmp[3684]*kernel[6]+tmp[3685]*kernel[7]+tmp[3686]*kernel[8];
				ans[3586]<=tmp[3485]*kernel[0]+tmp[3486]*kernel[1]+tmp[3487]*kernel[2]+tmp[3585]*kernel[3]+tmp[3586]*kernel[4]+tmp[3587]*kernel[5]+tmp[3685]*kernel[6]+tmp[3686]*kernel[7]+tmp[3687]*kernel[8];
				ans[3587]<=tmp[3486]*kernel[0]+tmp[3487]*kernel[1]+tmp[3488]*kernel[2]+tmp[3586]*kernel[3]+tmp[3587]*kernel[4]+tmp[3588]*kernel[5]+tmp[3686]*kernel[6]+tmp[3687]*kernel[7]+tmp[3688]*kernel[8];
				ans[3588]<=tmp[3487]*kernel[0]+tmp[3488]*kernel[1]+tmp[3489]*kernel[2]+tmp[3587]*kernel[3]+tmp[3588]*kernel[4]+tmp[3589]*kernel[5]+tmp[3687]*kernel[6]+tmp[3688]*kernel[7]+tmp[3689]*kernel[8];
				ans[3589]<=tmp[3488]*kernel[0]+tmp[3489]*kernel[1]+tmp[3490]*kernel[2]+tmp[3588]*kernel[3]+tmp[3589]*kernel[4]+tmp[3590]*kernel[5]+tmp[3688]*kernel[6]+tmp[3689]*kernel[7]+tmp[3690]*kernel[8];
				ans[3590]<=tmp[3489]*kernel[0]+tmp[3490]*kernel[1]+tmp[3491]*kernel[2]+tmp[3589]*kernel[3]+tmp[3590]*kernel[4]+tmp[3591]*kernel[5]+tmp[3689]*kernel[6]+tmp[3690]*kernel[7]+tmp[3691]*kernel[8];
				ans[3591]<=tmp[3490]*kernel[0]+tmp[3491]*kernel[1]+tmp[3492]*kernel[2]+tmp[3590]*kernel[3]+tmp[3591]*kernel[4]+tmp[3592]*kernel[5]+tmp[3690]*kernel[6]+tmp[3691]*kernel[7]+tmp[3692]*kernel[8];
				ans[3592]<=tmp[3491]*kernel[0]+tmp[3492]*kernel[1]+tmp[3493]*kernel[2]+tmp[3591]*kernel[3]+tmp[3592]*kernel[4]+tmp[3593]*kernel[5]+tmp[3691]*kernel[6]+tmp[3692]*kernel[7]+tmp[3693]*kernel[8];
				ans[3593]<=tmp[3492]*kernel[0]+tmp[3493]*kernel[1]+tmp[3494]*kernel[2]+tmp[3592]*kernel[3]+tmp[3593]*kernel[4]+tmp[3594]*kernel[5]+tmp[3692]*kernel[6]+tmp[3693]*kernel[7]+tmp[3694]*kernel[8];
				ans[3594]<=tmp[3493]*kernel[0]+tmp[3494]*kernel[1]+tmp[3495]*kernel[2]+tmp[3593]*kernel[3]+tmp[3594]*kernel[4]+tmp[3595]*kernel[5]+tmp[3693]*kernel[6]+tmp[3694]*kernel[7]+tmp[3695]*kernel[8];
				ans[3595]<=tmp[3494]*kernel[0]+tmp[3495]*kernel[1]+tmp[3496]*kernel[2]+tmp[3594]*kernel[3]+tmp[3595]*kernel[4]+tmp[3596]*kernel[5]+tmp[3694]*kernel[6]+tmp[3695]*kernel[7]+tmp[3696]*kernel[8];
				ans[3596]<=tmp[3495]*kernel[0]+tmp[3496]*kernel[1]+tmp[3497]*kernel[2]+tmp[3595]*kernel[3]+tmp[3596]*kernel[4]+tmp[3597]*kernel[5]+tmp[3695]*kernel[6]+tmp[3696]*kernel[7]+tmp[3697]*kernel[8];
				ans[3597]<=tmp[3496]*kernel[0]+tmp[3497]*kernel[1]+tmp[3498]*kernel[2]+tmp[3596]*kernel[3]+tmp[3597]*kernel[4]+tmp[3598]*kernel[5]+tmp[3696]*kernel[6]+tmp[3697]*kernel[7]+tmp[3698]*kernel[8];
				ans[3598]<=tmp[3497]*kernel[0]+tmp[3498]*kernel[1]+tmp[3499]*kernel[2]+tmp[3597]*kernel[3]+tmp[3598]*kernel[4]+tmp[3599]*kernel[5]+tmp[3697]*kernel[6]+tmp[3698]*kernel[7]+tmp[3699]*kernel[8];
				ans[3599]<=tmp[3498]*kernel[0]+tmp[3499]*kernel[1]+tmp[3598]*kernel[3]+tmp[3599]*kernel[4]+tmp[3698]*kernel[6]+tmp[3699]*kernel[7];
				ans[3600]<=tmp[3500]*kernel[1]+tmp[3501]*kernel[2]+tmp[3600]*kernel[4]+tmp[3601]*kernel[5]+tmp[3700]*kernel[7]+tmp[3701]*kernel[8];
				ans[3601]<=tmp[3500]*kernel[0]+tmp[3501]*kernel[1]+tmp[3502]*kernel[2]+tmp[3600]*kernel[3]+tmp[3601]*kernel[4]+tmp[3602]*kernel[5]+tmp[3700]*kernel[6]+tmp[3701]*kernel[7]+tmp[3702]*kernel[8];
				ans[3602]<=tmp[3501]*kernel[0]+tmp[3502]*kernel[1]+tmp[3503]*kernel[2]+tmp[3601]*kernel[3]+tmp[3602]*kernel[4]+tmp[3603]*kernel[5]+tmp[3701]*kernel[6]+tmp[3702]*kernel[7]+tmp[3703]*kernel[8];
				ans[3603]<=tmp[3502]*kernel[0]+tmp[3503]*kernel[1]+tmp[3504]*kernel[2]+tmp[3602]*kernel[3]+tmp[3603]*kernel[4]+tmp[3604]*kernel[5]+tmp[3702]*kernel[6]+tmp[3703]*kernel[7]+tmp[3704]*kernel[8];
				ans[3604]<=tmp[3503]*kernel[0]+tmp[3504]*kernel[1]+tmp[3505]*kernel[2]+tmp[3603]*kernel[3]+tmp[3604]*kernel[4]+tmp[3605]*kernel[5]+tmp[3703]*kernel[6]+tmp[3704]*kernel[7]+tmp[3705]*kernel[8];
				ans[3605]<=tmp[3504]*kernel[0]+tmp[3505]*kernel[1]+tmp[3506]*kernel[2]+tmp[3604]*kernel[3]+tmp[3605]*kernel[4]+tmp[3606]*kernel[5]+tmp[3704]*kernel[6]+tmp[3705]*kernel[7]+tmp[3706]*kernel[8];
				ans[3606]<=tmp[3505]*kernel[0]+tmp[3506]*kernel[1]+tmp[3507]*kernel[2]+tmp[3605]*kernel[3]+tmp[3606]*kernel[4]+tmp[3607]*kernel[5]+tmp[3705]*kernel[6]+tmp[3706]*kernel[7]+tmp[3707]*kernel[8];
				ans[3607]<=tmp[3506]*kernel[0]+tmp[3507]*kernel[1]+tmp[3508]*kernel[2]+tmp[3606]*kernel[3]+tmp[3607]*kernel[4]+tmp[3608]*kernel[5]+tmp[3706]*kernel[6]+tmp[3707]*kernel[7]+tmp[3708]*kernel[8];
				ans[3608]<=tmp[3507]*kernel[0]+tmp[3508]*kernel[1]+tmp[3509]*kernel[2]+tmp[3607]*kernel[3]+tmp[3608]*kernel[4]+tmp[3609]*kernel[5]+tmp[3707]*kernel[6]+tmp[3708]*kernel[7]+tmp[3709]*kernel[8];
				ans[3609]<=tmp[3508]*kernel[0]+tmp[3509]*kernel[1]+tmp[3510]*kernel[2]+tmp[3608]*kernel[3]+tmp[3609]*kernel[4]+tmp[3610]*kernel[5]+tmp[3708]*kernel[6]+tmp[3709]*kernel[7]+tmp[3710]*kernel[8];
				ans[3610]<=tmp[3509]*kernel[0]+tmp[3510]*kernel[1]+tmp[3511]*kernel[2]+tmp[3609]*kernel[3]+tmp[3610]*kernel[4]+tmp[3611]*kernel[5]+tmp[3709]*kernel[6]+tmp[3710]*kernel[7]+tmp[3711]*kernel[8];
				ans[3611]<=tmp[3510]*kernel[0]+tmp[3511]*kernel[1]+tmp[3512]*kernel[2]+tmp[3610]*kernel[3]+tmp[3611]*kernel[4]+tmp[3612]*kernel[5]+tmp[3710]*kernel[6]+tmp[3711]*kernel[7]+tmp[3712]*kernel[8];
				ans[3612]<=tmp[3511]*kernel[0]+tmp[3512]*kernel[1]+tmp[3513]*kernel[2]+tmp[3611]*kernel[3]+tmp[3612]*kernel[4]+tmp[3613]*kernel[5]+tmp[3711]*kernel[6]+tmp[3712]*kernel[7]+tmp[3713]*kernel[8];
				ans[3613]<=tmp[3512]*kernel[0]+tmp[3513]*kernel[1]+tmp[3514]*kernel[2]+tmp[3612]*kernel[3]+tmp[3613]*kernel[4]+tmp[3614]*kernel[5]+tmp[3712]*kernel[6]+tmp[3713]*kernel[7]+tmp[3714]*kernel[8];
				ans[3614]<=tmp[3513]*kernel[0]+tmp[3514]*kernel[1]+tmp[3515]*kernel[2]+tmp[3613]*kernel[3]+tmp[3614]*kernel[4]+tmp[3615]*kernel[5]+tmp[3713]*kernel[6]+tmp[3714]*kernel[7]+tmp[3715]*kernel[8];
				ans[3615]<=tmp[3514]*kernel[0]+tmp[3515]*kernel[1]+tmp[3516]*kernel[2]+tmp[3614]*kernel[3]+tmp[3615]*kernel[4]+tmp[3616]*kernel[5]+tmp[3714]*kernel[6]+tmp[3715]*kernel[7]+tmp[3716]*kernel[8];
				ans[3616]<=tmp[3515]*kernel[0]+tmp[3516]*kernel[1]+tmp[3517]*kernel[2]+tmp[3615]*kernel[3]+tmp[3616]*kernel[4]+tmp[3617]*kernel[5]+tmp[3715]*kernel[6]+tmp[3716]*kernel[7]+tmp[3717]*kernel[8];
				ans[3617]<=tmp[3516]*kernel[0]+tmp[3517]*kernel[1]+tmp[3518]*kernel[2]+tmp[3616]*kernel[3]+tmp[3617]*kernel[4]+tmp[3618]*kernel[5]+tmp[3716]*kernel[6]+tmp[3717]*kernel[7]+tmp[3718]*kernel[8];
				ans[3618]<=tmp[3517]*kernel[0]+tmp[3518]*kernel[1]+tmp[3519]*kernel[2]+tmp[3617]*kernel[3]+tmp[3618]*kernel[4]+tmp[3619]*kernel[5]+tmp[3717]*kernel[6]+tmp[3718]*kernel[7]+tmp[3719]*kernel[8];
				ans[3619]<=tmp[3518]*kernel[0]+tmp[3519]*kernel[1]+tmp[3520]*kernel[2]+tmp[3618]*kernel[3]+tmp[3619]*kernel[4]+tmp[3620]*kernel[5]+tmp[3718]*kernel[6]+tmp[3719]*kernel[7]+tmp[3720]*kernel[8];
				ans[3620]<=tmp[3519]*kernel[0]+tmp[3520]*kernel[1]+tmp[3521]*kernel[2]+tmp[3619]*kernel[3]+tmp[3620]*kernel[4]+tmp[3621]*kernel[5]+tmp[3719]*kernel[6]+tmp[3720]*kernel[7]+tmp[3721]*kernel[8];
				ans[3621]<=tmp[3520]*kernel[0]+tmp[3521]*kernel[1]+tmp[3522]*kernel[2]+tmp[3620]*kernel[3]+tmp[3621]*kernel[4]+tmp[3622]*kernel[5]+tmp[3720]*kernel[6]+tmp[3721]*kernel[7]+tmp[3722]*kernel[8];
				ans[3622]<=tmp[3521]*kernel[0]+tmp[3522]*kernel[1]+tmp[3523]*kernel[2]+tmp[3621]*kernel[3]+tmp[3622]*kernel[4]+tmp[3623]*kernel[5]+tmp[3721]*kernel[6]+tmp[3722]*kernel[7]+tmp[3723]*kernel[8];
				ans[3623]<=tmp[3522]*kernel[0]+tmp[3523]*kernel[1]+tmp[3524]*kernel[2]+tmp[3622]*kernel[3]+tmp[3623]*kernel[4]+tmp[3624]*kernel[5]+tmp[3722]*kernel[6]+tmp[3723]*kernel[7]+tmp[3724]*kernel[8];
				ans[3624]<=tmp[3523]*kernel[0]+tmp[3524]*kernel[1]+tmp[3525]*kernel[2]+tmp[3623]*kernel[3]+tmp[3624]*kernel[4]+tmp[3625]*kernel[5]+tmp[3723]*kernel[6]+tmp[3724]*kernel[7]+tmp[3725]*kernel[8];
				ans[3625]<=tmp[3524]*kernel[0]+tmp[3525]*kernel[1]+tmp[3526]*kernel[2]+tmp[3624]*kernel[3]+tmp[3625]*kernel[4]+tmp[3626]*kernel[5]+tmp[3724]*kernel[6]+tmp[3725]*kernel[7]+tmp[3726]*kernel[8];
				ans[3626]<=tmp[3525]*kernel[0]+tmp[3526]*kernel[1]+tmp[3527]*kernel[2]+tmp[3625]*kernel[3]+tmp[3626]*kernel[4]+tmp[3627]*kernel[5]+tmp[3725]*kernel[6]+tmp[3726]*kernel[7]+tmp[3727]*kernel[8];
				ans[3627]<=tmp[3526]*kernel[0]+tmp[3527]*kernel[1]+tmp[3528]*kernel[2]+tmp[3626]*kernel[3]+tmp[3627]*kernel[4]+tmp[3628]*kernel[5]+tmp[3726]*kernel[6]+tmp[3727]*kernel[7]+tmp[3728]*kernel[8];
				ans[3628]<=tmp[3527]*kernel[0]+tmp[3528]*kernel[1]+tmp[3529]*kernel[2]+tmp[3627]*kernel[3]+tmp[3628]*kernel[4]+tmp[3629]*kernel[5]+tmp[3727]*kernel[6]+tmp[3728]*kernel[7]+tmp[3729]*kernel[8];
				ans[3629]<=tmp[3528]*kernel[0]+tmp[3529]*kernel[1]+tmp[3530]*kernel[2]+tmp[3628]*kernel[3]+tmp[3629]*kernel[4]+tmp[3630]*kernel[5]+tmp[3728]*kernel[6]+tmp[3729]*kernel[7]+tmp[3730]*kernel[8];
				ans[3630]<=tmp[3529]*kernel[0]+tmp[3530]*kernel[1]+tmp[3531]*kernel[2]+tmp[3629]*kernel[3]+tmp[3630]*kernel[4]+tmp[3631]*kernel[5]+tmp[3729]*kernel[6]+tmp[3730]*kernel[7]+tmp[3731]*kernel[8];
				ans[3631]<=tmp[3530]*kernel[0]+tmp[3531]*kernel[1]+tmp[3532]*kernel[2]+tmp[3630]*kernel[3]+tmp[3631]*kernel[4]+tmp[3632]*kernel[5]+tmp[3730]*kernel[6]+tmp[3731]*kernel[7]+tmp[3732]*kernel[8];
				ans[3632]<=tmp[3531]*kernel[0]+tmp[3532]*kernel[1]+tmp[3533]*kernel[2]+tmp[3631]*kernel[3]+tmp[3632]*kernel[4]+tmp[3633]*kernel[5]+tmp[3731]*kernel[6]+tmp[3732]*kernel[7]+tmp[3733]*kernel[8];
				ans[3633]<=tmp[3532]*kernel[0]+tmp[3533]*kernel[1]+tmp[3534]*kernel[2]+tmp[3632]*kernel[3]+tmp[3633]*kernel[4]+tmp[3634]*kernel[5]+tmp[3732]*kernel[6]+tmp[3733]*kernel[7]+tmp[3734]*kernel[8];
				ans[3634]<=tmp[3533]*kernel[0]+tmp[3534]*kernel[1]+tmp[3535]*kernel[2]+tmp[3633]*kernel[3]+tmp[3634]*kernel[4]+tmp[3635]*kernel[5]+tmp[3733]*kernel[6]+tmp[3734]*kernel[7]+tmp[3735]*kernel[8];
				ans[3635]<=tmp[3534]*kernel[0]+tmp[3535]*kernel[1]+tmp[3536]*kernel[2]+tmp[3634]*kernel[3]+tmp[3635]*kernel[4]+tmp[3636]*kernel[5]+tmp[3734]*kernel[6]+tmp[3735]*kernel[7]+tmp[3736]*kernel[8];
				ans[3636]<=tmp[3535]*kernel[0]+tmp[3536]*kernel[1]+tmp[3537]*kernel[2]+tmp[3635]*kernel[3]+tmp[3636]*kernel[4]+tmp[3637]*kernel[5]+tmp[3735]*kernel[6]+tmp[3736]*kernel[7]+tmp[3737]*kernel[8];
				ans[3637]<=tmp[3536]*kernel[0]+tmp[3537]*kernel[1]+tmp[3538]*kernel[2]+tmp[3636]*kernel[3]+tmp[3637]*kernel[4]+tmp[3638]*kernel[5]+tmp[3736]*kernel[6]+tmp[3737]*kernel[7]+tmp[3738]*kernel[8];
				ans[3638]<=tmp[3537]*kernel[0]+tmp[3538]*kernel[1]+tmp[3539]*kernel[2]+tmp[3637]*kernel[3]+tmp[3638]*kernel[4]+tmp[3639]*kernel[5]+tmp[3737]*kernel[6]+tmp[3738]*kernel[7]+tmp[3739]*kernel[8];
				ans[3639]<=tmp[3538]*kernel[0]+tmp[3539]*kernel[1]+tmp[3540]*kernel[2]+tmp[3638]*kernel[3]+tmp[3639]*kernel[4]+tmp[3640]*kernel[5]+tmp[3738]*kernel[6]+tmp[3739]*kernel[7]+tmp[3740]*kernel[8];
				ans[3640]<=tmp[3539]*kernel[0]+tmp[3540]*kernel[1]+tmp[3541]*kernel[2]+tmp[3639]*kernel[3]+tmp[3640]*kernel[4]+tmp[3641]*kernel[5]+tmp[3739]*kernel[6]+tmp[3740]*kernel[7]+tmp[3741]*kernel[8];
				ans[3641]<=tmp[3540]*kernel[0]+tmp[3541]*kernel[1]+tmp[3542]*kernel[2]+tmp[3640]*kernel[3]+tmp[3641]*kernel[4]+tmp[3642]*kernel[5]+tmp[3740]*kernel[6]+tmp[3741]*kernel[7]+tmp[3742]*kernel[8];
				ans[3642]<=tmp[3541]*kernel[0]+tmp[3542]*kernel[1]+tmp[3543]*kernel[2]+tmp[3641]*kernel[3]+tmp[3642]*kernel[4]+tmp[3643]*kernel[5]+tmp[3741]*kernel[6]+tmp[3742]*kernel[7]+tmp[3743]*kernel[8];
				ans[3643]<=tmp[3542]*kernel[0]+tmp[3543]*kernel[1]+tmp[3544]*kernel[2]+tmp[3642]*kernel[3]+tmp[3643]*kernel[4]+tmp[3644]*kernel[5]+tmp[3742]*kernel[6]+tmp[3743]*kernel[7]+tmp[3744]*kernel[8];
				ans[3644]<=tmp[3543]*kernel[0]+tmp[3544]*kernel[1]+tmp[3545]*kernel[2]+tmp[3643]*kernel[3]+tmp[3644]*kernel[4]+tmp[3645]*kernel[5]+tmp[3743]*kernel[6]+tmp[3744]*kernel[7]+tmp[3745]*kernel[8];
				ans[3645]<=tmp[3544]*kernel[0]+tmp[3545]*kernel[1]+tmp[3546]*kernel[2]+tmp[3644]*kernel[3]+tmp[3645]*kernel[4]+tmp[3646]*kernel[5]+tmp[3744]*kernel[6]+tmp[3745]*kernel[7]+tmp[3746]*kernel[8];
				ans[3646]<=tmp[3545]*kernel[0]+tmp[3546]*kernel[1]+tmp[3547]*kernel[2]+tmp[3645]*kernel[3]+tmp[3646]*kernel[4]+tmp[3647]*kernel[5]+tmp[3745]*kernel[6]+tmp[3746]*kernel[7]+tmp[3747]*kernel[8];
				ans[3647]<=tmp[3546]*kernel[0]+tmp[3547]*kernel[1]+tmp[3548]*kernel[2]+tmp[3646]*kernel[3]+tmp[3647]*kernel[4]+tmp[3648]*kernel[5]+tmp[3746]*kernel[6]+tmp[3747]*kernel[7]+tmp[3748]*kernel[8];
				ans[3648]<=tmp[3547]*kernel[0]+tmp[3548]*kernel[1]+tmp[3549]*kernel[2]+tmp[3647]*kernel[3]+tmp[3648]*kernel[4]+tmp[3649]*kernel[5]+tmp[3747]*kernel[6]+tmp[3748]*kernel[7]+tmp[3749]*kernel[8];
				ans[3649]<=tmp[3548]*kernel[0]+tmp[3549]*kernel[1]+tmp[3550]*kernel[2]+tmp[3648]*kernel[3]+tmp[3649]*kernel[4]+tmp[3650]*kernel[5]+tmp[3748]*kernel[6]+tmp[3749]*kernel[7]+tmp[3750]*kernel[8];
				ans[3650]<=tmp[3549]*kernel[0]+tmp[3550]*kernel[1]+tmp[3551]*kernel[2]+tmp[3649]*kernel[3]+tmp[3650]*kernel[4]+tmp[3651]*kernel[5]+tmp[3749]*kernel[6]+tmp[3750]*kernel[7]+tmp[3751]*kernel[8];
				ans[3651]<=tmp[3550]*kernel[0]+tmp[3551]*kernel[1]+tmp[3552]*kernel[2]+tmp[3650]*kernel[3]+tmp[3651]*kernel[4]+tmp[3652]*kernel[5]+tmp[3750]*kernel[6]+tmp[3751]*kernel[7]+tmp[3752]*kernel[8];
				ans[3652]<=tmp[3551]*kernel[0]+tmp[3552]*kernel[1]+tmp[3553]*kernel[2]+tmp[3651]*kernel[3]+tmp[3652]*kernel[4]+tmp[3653]*kernel[5]+tmp[3751]*kernel[6]+tmp[3752]*kernel[7]+tmp[3753]*kernel[8];
				ans[3653]<=tmp[3552]*kernel[0]+tmp[3553]*kernel[1]+tmp[3554]*kernel[2]+tmp[3652]*kernel[3]+tmp[3653]*kernel[4]+tmp[3654]*kernel[5]+tmp[3752]*kernel[6]+tmp[3753]*kernel[7]+tmp[3754]*kernel[8];
				ans[3654]<=tmp[3553]*kernel[0]+tmp[3554]*kernel[1]+tmp[3555]*kernel[2]+tmp[3653]*kernel[3]+tmp[3654]*kernel[4]+tmp[3655]*kernel[5]+tmp[3753]*kernel[6]+tmp[3754]*kernel[7]+tmp[3755]*kernel[8];
				ans[3655]<=tmp[3554]*kernel[0]+tmp[3555]*kernel[1]+tmp[3556]*kernel[2]+tmp[3654]*kernel[3]+tmp[3655]*kernel[4]+tmp[3656]*kernel[5]+tmp[3754]*kernel[6]+tmp[3755]*kernel[7]+tmp[3756]*kernel[8];
				ans[3656]<=tmp[3555]*kernel[0]+tmp[3556]*kernel[1]+tmp[3557]*kernel[2]+tmp[3655]*kernel[3]+tmp[3656]*kernel[4]+tmp[3657]*kernel[5]+tmp[3755]*kernel[6]+tmp[3756]*kernel[7]+tmp[3757]*kernel[8];
				ans[3657]<=tmp[3556]*kernel[0]+tmp[3557]*kernel[1]+tmp[3558]*kernel[2]+tmp[3656]*kernel[3]+tmp[3657]*kernel[4]+tmp[3658]*kernel[5]+tmp[3756]*kernel[6]+tmp[3757]*kernel[7]+tmp[3758]*kernel[8];
				ans[3658]<=tmp[3557]*kernel[0]+tmp[3558]*kernel[1]+tmp[3559]*kernel[2]+tmp[3657]*kernel[3]+tmp[3658]*kernel[4]+tmp[3659]*kernel[5]+tmp[3757]*kernel[6]+tmp[3758]*kernel[7]+tmp[3759]*kernel[8];
				ans[3659]<=tmp[3558]*kernel[0]+tmp[3559]*kernel[1]+tmp[3560]*kernel[2]+tmp[3658]*kernel[3]+tmp[3659]*kernel[4]+tmp[3660]*kernel[5]+tmp[3758]*kernel[6]+tmp[3759]*kernel[7]+tmp[3760]*kernel[8];
				ans[3660]<=tmp[3559]*kernel[0]+tmp[3560]*kernel[1]+tmp[3561]*kernel[2]+tmp[3659]*kernel[3]+tmp[3660]*kernel[4]+tmp[3661]*kernel[5]+tmp[3759]*kernel[6]+tmp[3760]*kernel[7]+tmp[3761]*kernel[8];
				ans[3661]<=tmp[3560]*kernel[0]+tmp[3561]*kernel[1]+tmp[3562]*kernel[2]+tmp[3660]*kernel[3]+tmp[3661]*kernel[4]+tmp[3662]*kernel[5]+tmp[3760]*kernel[6]+tmp[3761]*kernel[7]+tmp[3762]*kernel[8];
				ans[3662]<=tmp[3561]*kernel[0]+tmp[3562]*kernel[1]+tmp[3563]*kernel[2]+tmp[3661]*kernel[3]+tmp[3662]*kernel[4]+tmp[3663]*kernel[5]+tmp[3761]*kernel[6]+tmp[3762]*kernel[7]+tmp[3763]*kernel[8];
				ans[3663]<=tmp[3562]*kernel[0]+tmp[3563]*kernel[1]+tmp[3564]*kernel[2]+tmp[3662]*kernel[3]+tmp[3663]*kernel[4]+tmp[3664]*kernel[5]+tmp[3762]*kernel[6]+tmp[3763]*kernel[7]+tmp[3764]*kernel[8];
				ans[3664]<=tmp[3563]*kernel[0]+tmp[3564]*kernel[1]+tmp[3565]*kernel[2]+tmp[3663]*kernel[3]+tmp[3664]*kernel[4]+tmp[3665]*kernel[5]+tmp[3763]*kernel[6]+tmp[3764]*kernel[7]+tmp[3765]*kernel[8];
				ans[3665]<=tmp[3564]*kernel[0]+tmp[3565]*kernel[1]+tmp[3566]*kernel[2]+tmp[3664]*kernel[3]+tmp[3665]*kernel[4]+tmp[3666]*kernel[5]+tmp[3764]*kernel[6]+tmp[3765]*kernel[7]+tmp[3766]*kernel[8];
				ans[3666]<=tmp[3565]*kernel[0]+tmp[3566]*kernel[1]+tmp[3567]*kernel[2]+tmp[3665]*kernel[3]+tmp[3666]*kernel[4]+tmp[3667]*kernel[5]+tmp[3765]*kernel[6]+tmp[3766]*kernel[7]+tmp[3767]*kernel[8];
				ans[3667]<=tmp[3566]*kernel[0]+tmp[3567]*kernel[1]+tmp[3568]*kernel[2]+tmp[3666]*kernel[3]+tmp[3667]*kernel[4]+tmp[3668]*kernel[5]+tmp[3766]*kernel[6]+tmp[3767]*kernel[7]+tmp[3768]*kernel[8];
				ans[3668]<=tmp[3567]*kernel[0]+tmp[3568]*kernel[1]+tmp[3569]*kernel[2]+tmp[3667]*kernel[3]+tmp[3668]*kernel[4]+tmp[3669]*kernel[5]+tmp[3767]*kernel[6]+tmp[3768]*kernel[7]+tmp[3769]*kernel[8];
				ans[3669]<=tmp[3568]*kernel[0]+tmp[3569]*kernel[1]+tmp[3570]*kernel[2]+tmp[3668]*kernel[3]+tmp[3669]*kernel[4]+tmp[3670]*kernel[5]+tmp[3768]*kernel[6]+tmp[3769]*kernel[7]+tmp[3770]*kernel[8];
				ans[3670]<=tmp[3569]*kernel[0]+tmp[3570]*kernel[1]+tmp[3571]*kernel[2]+tmp[3669]*kernel[3]+tmp[3670]*kernel[4]+tmp[3671]*kernel[5]+tmp[3769]*kernel[6]+tmp[3770]*kernel[7]+tmp[3771]*kernel[8];
				ans[3671]<=tmp[3570]*kernel[0]+tmp[3571]*kernel[1]+tmp[3572]*kernel[2]+tmp[3670]*kernel[3]+tmp[3671]*kernel[4]+tmp[3672]*kernel[5]+tmp[3770]*kernel[6]+tmp[3771]*kernel[7]+tmp[3772]*kernel[8];
				ans[3672]<=tmp[3571]*kernel[0]+tmp[3572]*kernel[1]+tmp[3573]*kernel[2]+tmp[3671]*kernel[3]+tmp[3672]*kernel[4]+tmp[3673]*kernel[5]+tmp[3771]*kernel[6]+tmp[3772]*kernel[7]+tmp[3773]*kernel[8];
				ans[3673]<=tmp[3572]*kernel[0]+tmp[3573]*kernel[1]+tmp[3574]*kernel[2]+tmp[3672]*kernel[3]+tmp[3673]*kernel[4]+tmp[3674]*kernel[5]+tmp[3772]*kernel[6]+tmp[3773]*kernel[7]+tmp[3774]*kernel[8];
				ans[3674]<=tmp[3573]*kernel[0]+tmp[3574]*kernel[1]+tmp[3575]*kernel[2]+tmp[3673]*kernel[3]+tmp[3674]*kernel[4]+tmp[3675]*kernel[5]+tmp[3773]*kernel[6]+tmp[3774]*kernel[7]+tmp[3775]*kernel[8];
				ans[3675]<=tmp[3574]*kernel[0]+tmp[3575]*kernel[1]+tmp[3576]*kernel[2]+tmp[3674]*kernel[3]+tmp[3675]*kernel[4]+tmp[3676]*kernel[5]+tmp[3774]*kernel[6]+tmp[3775]*kernel[7]+tmp[3776]*kernel[8];
				ans[3676]<=tmp[3575]*kernel[0]+tmp[3576]*kernel[1]+tmp[3577]*kernel[2]+tmp[3675]*kernel[3]+tmp[3676]*kernel[4]+tmp[3677]*kernel[5]+tmp[3775]*kernel[6]+tmp[3776]*kernel[7]+tmp[3777]*kernel[8];
				ans[3677]<=tmp[3576]*kernel[0]+tmp[3577]*kernel[1]+tmp[3578]*kernel[2]+tmp[3676]*kernel[3]+tmp[3677]*kernel[4]+tmp[3678]*kernel[5]+tmp[3776]*kernel[6]+tmp[3777]*kernel[7]+tmp[3778]*kernel[8];
				ans[3678]<=tmp[3577]*kernel[0]+tmp[3578]*kernel[1]+tmp[3579]*kernel[2]+tmp[3677]*kernel[3]+tmp[3678]*kernel[4]+tmp[3679]*kernel[5]+tmp[3777]*kernel[6]+tmp[3778]*kernel[7]+tmp[3779]*kernel[8];
				ans[3679]<=tmp[3578]*kernel[0]+tmp[3579]*kernel[1]+tmp[3580]*kernel[2]+tmp[3678]*kernel[3]+tmp[3679]*kernel[4]+tmp[3680]*kernel[5]+tmp[3778]*kernel[6]+tmp[3779]*kernel[7]+tmp[3780]*kernel[8];
				ans[3680]<=tmp[3579]*kernel[0]+tmp[3580]*kernel[1]+tmp[3581]*kernel[2]+tmp[3679]*kernel[3]+tmp[3680]*kernel[4]+tmp[3681]*kernel[5]+tmp[3779]*kernel[6]+tmp[3780]*kernel[7]+tmp[3781]*kernel[8];
				ans[3681]<=tmp[3580]*kernel[0]+tmp[3581]*kernel[1]+tmp[3582]*kernel[2]+tmp[3680]*kernel[3]+tmp[3681]*kernel[4]+tmp[3682]*kernel[5]+tmp[3780]*kernel[6]+tmp[3781]*kernel[7]+tmp[3782]*kernel[8];
				ans[3682]<=tmp[3581]*kernel[0]+tmp[3582]*kernel[1]+tmp[3583]*kernel[2]+tmp[3681]*kernel[3]+tmp[3682]*kernel[4]+tmp[3683]*kernel[5]+tmp[3781]*kernel[6]+tmp[3782]*kernel[7]+tmp[3783]*kernel[8];
				ans[3683]<=tmp[3582]*kernel[0]+tmp[3583]*kernel[1]+tmp[3584]*kernel[2]+tmp[3682]*kernel[3]+tmp[3683]*kernel[4]+tmp[3684]*kernel[5]+tmp[3782]*kernel[6]+tmp[3783]*kernel[7]+tmp[3784]*kernel[8];
				ans[3684]<=tmp[3583]*kernel[0]+tmp[3584]*kernel[1]+tmp[3585]*kernel[2]+tmp[3683]*kernel[3]+tmp[3684]*kernel[4]+tmp[3685]*kernel[5]+tmp[3783]*kernel[6]+tmp[3784]*kernel[7]+tmp[3785]*kernel[8];
				ans[3685]<=tmp[3584]*kernel[0]+tmp[3585]*kernel[1]+tmp[3586]*kernel[2]+tmp[3684]*kernel[3]+tmp[3685]*kernel[4]+tmp[3686]*kernel[5]+tmp[3784]*kernel[6]+tmp[3785]*kernel[7]+tmp[3786]*kernel[8];
				ans[3686]<=tmp[3585]*kernel[0]+tmp[3586]*kernel[1]+tmp[3587]*kernel[2]+tmp[3685]*kernel[3]+tmp[3686]*kernel[4]+tmp[3687]*kernel[5]+tmp[3785]*kernel[6]+tmp[3786]*kernel[7]+tmp[3787]*kernel[8];
				ans[3687]<=tmp[3586]*kernel[0]+tmp[3587]*kernel[1]+tmp[3588]*kernel[2]+tmp[3686]*kernel[3]+tmp[3687]*kernel[4]+tmp[3688]*kernel[5]+tmp[3786]*kernel[6]+tmp[3787]*kernel[7]+tmp[3788]*kernel[8];
				ans[3688]<=tmp[3587]*kernel[0]+tmp[3588]*kernel[1]+tmp[3589]*kernel[2]+tmp[3687]*kernel[3]+tmp[3688]*kernel[4]+tmp[3689]*kernel[5]+tmp[3787]*kernel[6]+tmp[3788]*kernel[7]+tmp[3789]*kernel[8];
				ans[3689]<=tmp[3588]*kernel[0]+tmp[3589]*kernel[1]+tmp[3590]*kernel[2]+tmp[3688]*kernel[3]+tmp[3689]*kernel[4]+tmp[3690]*kernel[5]+tmp[3788]*kernel[6]+tmp[3789]*kernel[7]+tmp[3790]*kernel[8];
				ans[3690]<=tmp[3589]*kernel[0]+tmp[3590]*kernel[1]+tmp[3591]*kernel[2]+tmp[3689]*kernel[3]+tmp[3690]*kernel[4]+tmp[3691]*kernel[5]+tmp[3789]*kernel[6]+tmp[3790]*kernel[7]+tmp[3791]*kernel[8];
				ans[3691]<=tmp[3590]*kernel[0]+tmp[3591]*kernel[1]+tmp[3592]*kernel[2]+tmp[3690]*kernel[3]+tmp[3691]*kernel[4]+tmp[3692]*kernel[5]+tmp[3790]*kernel[6]+tmp[3791]*kernel[7]+tmp[3792]*kernel[8];
				ans[3692]<=tmp[3591]*kernel[0]+tmp[3592]*kernel[1]+tmp[3593]*kernel[2]+tmp[3691]*kernel[3]+tmp[3692]*kernel[4]+tmp[3693]*kernel[5]+tmp[3791]*kernel[6]+tmp[3792]*kernel[7]+tmp[3793]*kernel[8];
				ans[3693]<=tmp[3592]*kernel[0]+tmp[3593]*kernel[1]+tmp[3594]*kernel[2]+tmp[3692]*kernel[3]+tmp[3693]*kernel[4]+tmp[3694]*kernel[5]+tmp[3792]*kernel[6]+tmp[3793]*kernel[7]+tmp[3794]*kernel[8];
				ans[3694]<=tmp[3593]*kernel[0]+tmp[3594]*kernel[1]+tmp[3595]*kernel[2]+tmp[3693]*kernel[3]+tmp[3694]*kernel[4]+tmp[3695]*kernel[5]+tmp[3793]*kernel[6]+tmp[3794]*kernel[7]+tmp[3795]*kernel[8];
				ans[3695]<=tmp[3594]*kernel[0]+tmp[3595]*kernel[1]+tmp[3596]*kernel[2]+tmp[3694]*kernel[3]+tmp[3695]*kernel[4]+tmp[3696]*kernel[5]+tmp[3794]*kernel[6]+tmp[3795]*kernel[7]+tmp[3796]*kernel[8];
				ans[3696]<=tmp[3595]*kernel[0]+tmp[3596]*kernel[1]+tmp[3597]*kernel[2]+tmp[3695]*kernel[3]+tmp[3696]*kernel[4]+tmp[3697]*kernel[5]+tmp[3795]*kernel[6]+tmp[3796]*kernel[7]+tmp[3797]*kernel[8];
				ans[3697]<=tmp[3596]*kernel[0]+tmp[3597]*kernel[1]+tmp[3598]*kernel[2]+tmp[3696]*kernel[3]+tmp[3697]*kernel[4]+tmp[3698]*kernel[5]+tmp[3796]*kernel[6]+tmp[3797]*kernel[7]+tmp[3798]*kernel[8];
				ans[3698]<=tmp[3597]*kernel[0]+tmp[3598]*kernel[1]+tmp[3599]*kernel[2]+tmp[3697]*kernel[3]+tmp[3698]*kernel[4]+tmp[3699]*kernel[5]+tmp[3797]*kernel[6]+tmp[3798]*kernel[7]+tmp[3799]*kernel[8];
				ans[3699]<=tmp[3598]*kernel[0]+tmp[3599]*kernel[1]+tmp[3698]*kernel[3]+tmp[3699]*kernel[4]+tmp[3798]*kernel[6]+tmp[3799]*kernel[7];
				ans[3700]<=tmp[3600]*kernel[1]+tmp[3601]*kernel[2]+tmp[3700]*kernel[4]+tmp[3701]*kernel[5]+tmp[3800]*kernel[7]+tmp[3801]*kernel[8];
				ans[3701]<=tmp[3600]*kernel[0]+tmp[3601]*kernel[1]+tmp[3602]*kernel[2]+tmp[3700]*kernel[3]+tmp[3701]*kernel[4]+tmp[3702]*kernel[5]+tmp[3800]*kernel[6]+tmp[3801]*kernel[7]+tmp[3802]*kernel[8];
				ans[3702]<=tmp[3601]*kernel[0]+tmp[3602]*kernel[1]+tmp[3603]*kernel[2]+tmp[3701]*kernel[3]+tmp[3702]*kernel[4]+tmp[3703]*kernel[5]+tmp[3801]*kernel[6]+tmp[3802]*kernel[7]+tmp[3803]*kernel[8];
				ans[3703]<=tmp[3602]*kernel[0]+tmp[3603]*kernel[1]+tmp[3604]*kernel[2]+tmp[3702]*kernel[3]+tmp[3703]*kernel[4]+tmp[3704]*kernel[5]+tmp[3802]*kernel[6]+tmp[3803]*kernel[7]+tmp[3804]*kernel[8];
				ans[3704]<=tmp[3603]*kernel[0]+tmp[3604]*kernel[1]+tmp[3605]*kernel[2]+tmp[3703]*kernel[3]+tmp[3704]*kernel[4]+tmp[3705]*kernel[5]+tmp[3803]*kernel[6]+tmp[3804]*kernel[7]+tmp[3805]*kernel[8];
				ans[3705]<=tmp[3604]*kernel[0]+tmp[3605]*kernel[1]+tmp[3606]*kernel[2]+tmp[3704]*kernel[3]+tmp[3705]*kernel[4]+tmp[3706]*kernel[5]+tmp[3804]*kernel[6]+tmp[3805]*kernel[7]+tmp[3806]*kernel[8];
				ans[3706]<=tmp[3605]*kernel[0]+tmp[3606]*kernel[1]+tmp[3607]*kernel[2]+tmp[3705]*kernel[3]+tmp[3706]*kernel[4]+tmp[3707]*kernel[5]+tmp[3805]*kernel[6]+tmp[3806]*kernel[7]+tmp[3807]*kernel[8];
				ans[3707]<=tmp[3606]*kernel[0]+tmp[3607]*kernel[1]+tmp[3608]*kernel[2]+tmp[3706]*kernel[3]+tmp[3707]*kernel[4]+tmp[3708]*kernel[5]+tmp[3806]*kernel[6]+tmp[3807]*kernel[7]+tmp[3808]*kernel[8];
				ans[3708]<=tmp[3607]*kernel[0]+tmp[3608]*kernel[1]+tmp[3609]*kernel[2]+tmp[3707]*kernel[3]+tmp[3708]*kernel[4]+tmp[3709]*kernel[5]+tmp[3807]*kernel[6]+tmp[3808]*kernel[7]+tmp[3809]*kernel[8];
				ans[3709]<=tmp[3608]*kernel[0]+tmp[3609]*kernel[1]+tmp[3610]*kernel[2]+tmp[3708]*kernel[3]+tmp[3709]*kernel[4]+tmp[3710]*kernel[5]+tmp[3808]*kernel[6]+tmp[3809]*kernel[7]+tmp[3810]*kernel[8];
				ans[3710]<=tmp[3609]*kernel[0]+tmp[3610]*kernel[1]+tmp[3611]*kernel[2]+tmp[3709]*kernel[3]+tmp[3710]*kernel[4]+tmp[3711]*kernel[5]+tmp[3809]*kernel[6]+tmp[3810]*kernel[7]+tmp[3811]*kernel[8];
				ans[3711]<=tmp[3610]*kernel[0]+tmp[3611]*kernel[1]+tmp[3612]*kernel[2]+tmp[3710]*kernel[3]+tmp[3711]*kernel[4]+tmp[3712]*kernel[5]+tmp[3810]*kernel[6]+tmp[3811]*kernel[7]+tmp[3812]*kernel[8];
				ans[3712]<=tmp[3611]*kernel[0]+tmp[3612]*kernel[1]+tmp[3613]*kernel[2]+tmp[3711]*kernel[3]+tmp[3712]*kernel[4]+tmp[3713]*kernel[5]+tmp[3811]*kernel[6]+tmp[3812]*kernel[7]+tmp[3813]*kernel[8];
				ans[3713]<=tmp[3612]*kernel[0]+tmp[3613]*kernel[1]+tmp[3614]*kernel[2]+tmp[3712]*kernel[3]+tmp[3713]*kernel[4]+tmp[3714]*kernel[5]+tmp[3812]*kernel[6]+tmp[3813]*kernel[7]+tmp[3814]*kernel[8];
				ans[3714]<=tmp[3613]*kernel[0]+tmp[3614]*kernel[1]+tmp[3615]*kernel[2]+tmp[3713]*kernel[3]+tmp[3714]*kernel[4]+tmp[3715]*kernel[5]+tmp[3813]*kernel[6]+tmp[3814]*kernel[7]+tmp[3815]*kernel[8];
				ans[3715]<=tmp[3614]*kernel[0]+tmp[3615]*kernel[1]+tmp[3616]*kernel[2]+tmp[3714]*kernel[3]+tmp[3715]*kernel[4]+tmp[3716]*kernel[5]+tmp[3814]*kernel[6]+tmp[3815]*kernel[7]+tmp[3816]*kernel[8];
				ans[3716]<=tmp[3615]*kernel[0]+tmp[3616]*kernel[1]+tmp[3617]*kernel[2]+tmp[3715]*kernel[3]+tmp[3716]*kernel[4]+tmp[3717]*kernel[5]+tmp[3815]*kernel[6]+tmp[3816]*kernel[7]+tmp[3817]*kernel[8];
				ans[3717]<=tmp[3616]*kernel[0]+tmp[3617]*kernel[1]+tmp[3618]*kernel[2]+tmp[3716]*kernel[3]+tmp[3717]*kernel[4]+tmp[3718]*kernel[5]+tmp[3816]*kernel[6]+tmp[3817]*kernel[7]+tmp[3818]*kernel[8];
				ans[3718]<=tmp[3617]*kernel[0]+tmp[3618]*kernel[1]+tmp[3619]*kernel[2]+tmp[3717]*kernel[3]+tmp[3718]*kernel[4]+tmp[3719]*kernel[5]+tmp[3817]*kernel[6]+tmp[3818]*kernel[7]+tmp[3819]*kernel[8];
				ans[3719]<=tmp[3618]*kernel[0]+tmp[3619]*kernel[1]+tmp[3620]*kernel[2]+tmp[3718]*kernel[3]+tmp[3719]*kernel[4]+tmp[3720]*kernel[5]+tmp[3818]*kernel[6]+tmp[3819]*kernel[7]+tmp[3820]*kernel[8];
				ans[3720]<=tmp[3619]*kernel[0]+tmp[3620]*kernel[1]+tmp[3621]*kernel[2]+tmp[3719]*kernel[3]+tmp[3720]*kernel[4]+tmp[3721]*kernel[5]+tmp[3819]*kernel[6]+tmp[3820]*kernel[7]+tmp[3821]*kernel[8];
				ans[3721]<=tmp[3620]*kernel[0]+tmp[3621]*kernel[1]+tmp[3622]*kernel[2]+tmp[3720]*kernel[3]+tmp[3721]*kernel[4]+tmp[3722]*kernel[5]+tmp[3820]*kernel[6]+tmp[3821]*kernel[7]+tmp[3822]*kernel[8];
				ans[3722]<=tmp[3621]*kernel[0]+tmp[3622]*kernel[1]+tmp[3623]*kernel[2]+tmp[3721]*kernel[3]+tmp[3722]*kernel[4]+tmp[3723]*kernel[5]+tmp[3821]*kernel[6]+tmp[3822]*kernel[7]+tmp[3823]*kernel[8];
				ans[3723]<=tmp[3622]*kernel[0]+tmp[3623]*kernel[1]+tmp[3624]*kernel[2]+tmp[3722]*kernel[3]+tmp[3723]*kernel[4]+tmp[3724]*kernel[5]+tmp[3822]*kernel[6]+tmp[3823]*kernel[7]+tmp[3824]*kernel[8];
				ans[3724]<=tmp[3623]*kernel[0]+tmp[3624]*kernel[1]+tmp[3625]*kernel[2]+tmp[3723]*kernel[3]+tmp[3724]*kernel[4]+tmp[3725]*kernel[5]+tmp[3823]*kernel[6]+tmp[3824]*kernel[7]+tmp[3825]*kernel[8];
				ans[3725]<=tmp[3624]*kernel[0]+tmp[3625]*kernel[1]+tmp[3626]*kernel[2]+tmp[3724]*kernel[3]+tmp[3725]*kernel[4]+tmp[3726]*kernel[5]+tmp[3824]*kernel[6]+tmp[3825]*kernel[7]+tmp[3826]*kernel[8];
				ans[3726]<=tmp[3625]*kernel[0]+tmp[3626]*kernel[1]+tmp[3627]*kernel[2]+tmp[3725]*kernel[3]+tmp[3726]*kernel[4]+tmp[3727]*kernel[5]+tmp[3825]*kernel[6]+tmp[3826]*kernel[7]+tmp[3827]*kernel[8];
				ans[3727]<=tmp[3626]*kernel[0]+tmp[3627]*kernel[1]+tmp[3628]*kernel[2]+tmp[3726]*kernel[3]+tmp[3727]*kernel[4]+tmp[3728]*kernel[5]+tmp[3826]*kernel[6]+tmp[3827]*kernel[7]+tmp[3828]*kernel[8];
				ans[3728]<=tmp[3627]*kernel[0]+tmp[3628]*kernel[1]+tmp[3629]*kernel[2]+tmp[3727]*kernel[3]+tmp[3728]*kernel[4]+tmp[3729]*kernel[5]+tmp[3827]*kernel[6]+tmp[3828]*kernel[7]+tmp[3829]*kernel[8];
				ans[3729]<=tmp[3628]*kernel[0]+tmp[3629]*kernel[1]+tmp[3630]*kernel[2]+tmp[3728]*kernel[3]+tmp[3729]*kernel[4]+tmp[3730]*kernel[5]+tmp[3828]*kernel[6]+tmp[3829]*kernel[7]+tmp[3830]*kernel[8];
				ans[3730]<=tmp[3629]*kernel[0]+tmp[3630]*kernel[1]+tmp[3631]*kernel[2]+tmp[3729]*kernel[3]+tmp[3730]*kernel[4]+tmp[3731]*kernel[5]+tmp[3829]*kernel[6]+tmp[3830]*kernel[7]+tmp[3831]*kernel[8];
				ans[3731]<=tmp[3630]*kernel[0]+tmp[3631]*kernel[1]+tmp[3632]*kernel[2]+tmp[3730]*kernel[3]+tmp[3731]*kernel[4]+tmp[3732]*kernel[5]+tmp[3830]*kernel[6]+tmp[3831]*kernel[7]+tmp[3832]*kernel[8];
				ans[3732]<=tmp[3631]*kernel[0]+tmp[3632]*kernel[1]+tmp[3633]*kernel[2]+tmp[3731]*kernel[3]+tmp[3732]*kernel[4]+tmp[3733]*kernel[5]+tmp[3831]*kernel[6]+tmp[3832]*kernel[7]+tmp[3833]*kernel[8];
				ans[3733]<=tmp[3632]*kernel[0]+tmp[3633]*kernel[1]+tmp[3634]*kernel[2]+tmp[3732]*kernel[3]+tmp[3733]*kernel[4]+tmp[3734]*kernel[5]+tmp[3832]*kernel[6]+tmp[3833]*kernel[7]+tmp[3834]*kernel[8];
				ans[3734]<=tmp[3633]*kernel[0]+tmp[3634]*kernel[1]+tmp[3635]*kernel[2]+tmp[3733]*kernel[3]+tmp[3734]*kernel[4]+tmp[3735]*kernel[5]+tmp[3833]*kernel[6]+tmp[3834]*kernel[7]+tmp[3835]*kernel[8];
				ans[3735]<=tmp[3634]*kernel[0]+tmp[3635]*kernel[1]+tmp[3636]*kernel[2]+tmp[3734]*kernel[3]+tmp[3735]*kernel[4]+tmp[3736]*kernel[5]+tmp[3834]*kernel[6]+tmp[3835]*kernel[7]+tmp[3836]*kernel[8];
				ans[3736]<=tmp[3635]*kernel[0]+tmp[3636]*kernel[1]+tmp[3637]*kernel[2]+tmp[3735]*kernel[3]+tmp[3736]*kernel[4]+tmp[3737]*kernel[5]+tmp[3835]*kernel[6]+tmp[3836]*kernel[7]+tmp[3837]*kernel[8];
				ans[3737]<=tmp[3636]*kernel[0]+tmp[3637]*kernel[1]+tmp[3638]*kernel[2]+tmp[3736]*kernel[3]+tmp[3737]*kernel[4]+tmp[3738]*kernel[5]+tmp[3836]*kernel[6]+tmp[3837]*kernel[7]+tmp[3838]*kernel[8];
				ans[3738]<=tmp[3637]*kernel[0]+tmp[3638]*kernel[1]+tmp[3639]*kernel[2]+tmp[3737]*kernel[3]+tmp[3738]*kernel[4]+tmp[3739]*kernel[5]+tmp[3837]*kernel[6]+tmp[3838]*kernel[7]+tmp[3839]*kernel[8];
				ans[3739]<=tmp[3638]*kernel[0]+tmp[3639]*kernel[1]+tmp[3640]*kernel[2]+tmp[3738]*kernel[3]+tmp[3739]*kernel[4]+tmp[3740]*kernel[5]+tmp[3838]*kernel[6]+tmp[3839]*kernel[7]+tmp[3840]*kernel[8];
				ans[3740]<=tmp[3639]*kernel[0]+tmp[3640]*kernel[1]+tmp[3641]*kernel[2]+tmp[3739]*kernel[3]+tmp[3740]*kernel[4]+tmp[3741]*kernel[5]+tmp[3839]*kernel[6]+tmp[3840]*kernel[7]+tmp[3841]*kernel[8];
				ans[3741]<=tmp[3640]*kernel[0]+tmp[3641]*kernel[1]+tmp[3642]*kernel[2]+tmp[3740]*kernel[3]+tmp[3741]*kernel[4]+tmp[3742]*kernel[5]+tmp[3840]*kernel[6]+tmp[3841]*kernel[7]+tmp[3842]*kernel[8];
				ans[3742]<=tmp[3641]*kernel[0]+tmp[3642]*kernel[1]+tmp[3643]*kernel[2]+tmp[3741]*kernel[3]+tmp[3742]*kernel[4]+tmp[3743]*kernel[5]+tmp[3841]*kernel[6]+tmp[3842]*kernel[7]+tmp[3843]*kernel[8];
				ans[3743]<=tmp[3642]*kernel[0]+tmp[3643]*kernel[1]+tmp[3644]*kernel[2]+tmp[3742]*kernel[3]+tmp[3743]*kernel[4]+tmp[3744]*kernel[5]+tmp[3842]*kernel[6]+tmp[3843]*kernel[7]+tmp[3844]*kernel[8];
				ans[3744]<=tmp[3643]*kernel[0]+tmp[3644]*kernel[1]+tmp[3645]*kernel[2]+tmp[3743]*kernel[3]+tmp[3744]*kernel[4]+tmp[3745]*kernel[5]+tmp[3843]*kernel[6]+tmp[3844]*kernel[7]+tmp[3845]*kernel[8];
				ans[3745]<=tmp[3644]*kernel[0]+tmp[3645]*kernel[1]+tmp[3646]*kernel[2]+tmp[3744]*kernel[3]+tmp[3745]*kernel[4]+tmp[3746]*kernel[5]+tmp[3844]*kernel[6]+tmp[3845]*kernel[7]+tmp[3846]*kernel[8];
				ans[3746]<=tmp[3645]*kernel[0]+tmp[3646]*kernel[1]+tmp[3647]*kernel[2]+tmp[3745]*kernel[3]+tmp[3746]*kernel[4]+tmp[3747]*kernel[5]+tmp[3845]*kernel[6]+tmp[3846]*kernel[7]+tmp[3847]*kernel[8];
				ans[3747]<=tmp[3646]*kernel[0]+tmp[3647]*kernel[1]+tmp[3648]*kernel[2]+tmp[3746]*kernel[3]+tmp[3747]*kernel[4]+tmp[3748]*kernel[5]+tmp[3846]*kernel[6]+tmp[3847]*kernel[7]+tmp[3848]*kernel[8];
				ans[3748]<=tmp[3647]*kernel[0]+tmp[3648]*kernel[1]+tmp[3649]*kernel[2]+tmp[3747]*kernel[3]+tmp[3748]*kernel[4]+tmp[3749]*kernel[5]+tmp[3847]*kernel[6]+tmp[3848]*kernel[7]+tmp[3849]*kernel[8];
				ans[3749]<=tmp[3648]*kernel[0]+tmp[3649]*kernel[1]+tmp[3650]*kernel[2]+tmp[3748]*kernel[3]+tmp[3749]*kernel[4]+tmp[3750]*kernel[5]+tmp[3848]*kernel[6]+tmp[3849]*kernel[7]+tmp[3850]*kernel[8];
				ans[3750]<=tmp[3649]*kernel[0]+tmp[3650]*kernel[1]+tmp[3651]*kernel[2]+tmp[3749]*kernel[3]+tmp[3750]*kernel[4]+tmp[3751]*kernel[5]+tmp[3849]*kernel[6]+tmp[3850]*kernel[7]+tmp[3851]*kernel[8];
				ans[3751]<=tmp[3650]*kernel[0]+tmp[3651]*kernel[1]+tmp[3652]*kernel[2]+tmp[3750]*kernel[3]+tmp[3751]*kernel[4]+tmp[3752]*kernel[5]+tmp[3850]*kernel[6]+tmp[3851]*kernel[7]+tmp[3852]*kernel[8];
				ans[3752]<=tmp[3651]*kernel[0]+tmp[3652]*kernel[1]+tmp[3653]*kernel[2]+tmp[3751]*kernel[3]+tmp[3752]*kernel[4]+tmp[3753]*kernel[5]+tmp[3851]*kernel[6]+tmp[3852]*kernel[7]+tmp[3853]*kernel[8];
				ans[3753]<=tmp[3652]*kernel[0]+tmp[3653]*kernel[1]+tmp[3654]*kernel[2]+tmp[3752]*kernel[3]+tmp[3753]*kernel[4]+tmp[3754]*kernel[5]+tmp[3852]*kernel[6]+tmp[3853]*kernel[7]+tmp[3854]*kernel[8];
				ans[3754]<=tmp[3653]*kernel[0]+tmp[3654]*kernel[1]+tmp[3655]*kernel[2]+tmp[3753]*kernel[3]+tmp[3754]*kernel[4]+tmp[3755]*kernel[5]+tmp[3853]*kernel[6]+tmp[3854]*kernel[7]+tmp[3855]*kernel[8];
				ans[3755]<=tmp[3654]*kernel[0]+tmp[3655]*kernel[1]+tmp[3656]*kernel[2]+tmp[3754]*kernel[3]+tmp[3755]*kernel[4]+tmp[3756]*kernel[5]+tmp[3854]*kernel[6]+tmp[3855]*kernel[7]+tmp[3856]*kernel[8];
				ans[3756]<=tmp[3655]*kernel[0]+tmp[3656]*kernel[1]+tmp[3657]*kernel[2]+tmp[3755]*kernel[3]+tmp[3756]*kernel[4]+tmp[3757]*kernel[5]+tmp[3855]*kernel[6]+tmp[3856]*kernel[7]+tmp[3857]*kernel[8];
				ans[3757]<=tmp[3656]*kernel[0]+tmp[3657]*kernel[1]+tmp[3658]*kernel[2]+tmp[3756]*kernel[3]+tmp[3757]*kernel[4]+tmp[3758]*kernel[5]+tmp[3856]*kernel[6]+tmp[3857]*kernel[7]+tmp[3858]*kernel[8];
				ans[3758]<=tmp[3657]*kernel[0]+tmp[3658]*kernel[1]+tmp[3659]*kernel[2]+tmp[3757]*kernel[3]+tmp[3758]*kernel[4]+tmp[3759]*kernel[5]+tmp[3857]*kernel[6]+tmp[3858]*kernel[7]+tmp[3859]*kernel[8];
				ans[3759]<=tmp[3658]*kernel[0]+tmp[3659]*kernel[1]+tmp[3660]*kernel[2]+tmp[3758]*kernel[3]+tmp[3759]*kernel[4]+tmp[3760]*kernel[5]+tmp[3858]*kernel[6]+tmp[3859]*kernel[7]+tmp[3860]*kernel[8];
				ans[3760]<=tmp[3659]*kernel[0]+tmp[3660]*kernel[1]+tmp[3661]*kernel[2]+tmp[3759]*kernel[3]+tmp[3760]*kernel[4]+tmp[3761]*kernel[5]+tmp[3859]*kernel[6]+tmp[3860]*kernel[7]+tmp[3861]*kernel[8];
				ans[3761]<=tmp[3660]*kernel[0]+tmp[3661]*kernel[1]+tmp[3662]*kernel[2]+tmp[3760]*kernel[3]+tmp[3761]*kernel[4]+tmp[3762]*kernel[5]+tmp[3860]*kernel[6]+tmp[3861]*kernel[7]+tmp[3862]*kernel[8];
				ans[3762]<=tmp[3661]*kernel[0]+tmp[3662]*kernel[1]+tmp[3663]*kernel[2]+tmp[3761]*kernel[3]+tmp[3762]*kernel[4]+tmp[3763]*kernel[5]+tmp[3861]*kernel[6]+tmp[3862]*kernel[7]+tmp[3863]*kernel[8];
				ans[3763]<=tmp[3662]*kernel[0]+tmp[3663]*kernel[1]+tmp[3664]*kernel[2]+tmp[3762]*kernel[3]+tmp[3763]*kernel[4]+tmp[3764]*kernel[5]+tmp[3862]*kernel[6]+tmp[3863]*kernel[7]+tmp[3864]*kernel[8];
				ans[3764]<=tmp[3663]*kernel[0]+tmp[3664]*kernel[1]+tmp[3665]*kernel[2]+tmp[3763]*kernel[3]+tmp[3764]*kernel[4]+tmp[3765]*kernel[5]+tmp[3863]*kernel[6]+tmp[3864]*kernel[7]+tmp[3865]*kernel[8];
				ans[3765]<=tmp[3664]*kernel[0]+tmp[3665]*kernel[1]+tmp[3666]*kernel[2]+tmp[3764]*kernel[3]+tmp[3765]*kernel[4]+tmp[3766]*kernel[5]+tmp[3864]*kernel[6]+tmp[3865]*kernel[7]+tmp[3866]*kernel[8];
				ans[3766]<=tmp[3665]*kernel[0]+tmp[3666]*kernel[1]+tmp[3667]*kernel[2]+tmp[3765]*kernel[3]+tmp[3766]*kernel[4]+tmp[3767]*kernel[5]+tmp[3865]*kernel[6]+tmp[3866]*kernel[7]+tmp[3867]*kernel[8];
				ans[3767]<=tmp[3666]*kernel[0]+tmp[3667]*kernel[1]+tmp[3668]*kernel[2]+tmp[3766]*kernel[3]+tmp[3767]*kernel[4]+tmp[3768]*kernel[5]+tmp[3866]*kernel[6]+tmp[3867]*kernel[7]+tmp[3868]*kernel[8];
				ans[3768]<=tmp[3667]*kernel[0]+tmp[3668]*kernel[1]+tmp[3669]*kernel[2]+tmp[3767]*kernel[3]+tmp[3768]*kernel[4]+tmp[3769]*kernel[5]+tmp[3867]*kernel[6]+tmp[3868]*kernel[7]+tmp[3869]*kernel[8];
				ans[3769]<=tmp[3668]*kernel[0]+tmp[3669]*kernel[1]+tmp[3670]*kernel[2]+tmp[3768]*kernel[3]+tmp[3769]*kernel[4]+tmp[3770]*kernel[5]+tmp[3868]*kernel[6]+tmp[3869]*kernel[7]+tmp[3870]*kernel[8];
				ans[3770]<=tmp[3669]*kernel[0]+tmp[3670]*kernel[1]+tmp[3671]*kernel[2]+tmp[3769]*kernel[3]+tmp[3770]*kernel[4]+tmp[3771]*kernel[5]+tmp[3869]*kernel[6]+tmp[3870]*kernel[7]+tmp[3871]*kernel[8];
				ans[3771]<=tmp[3670]*kernel[0]+tmp[3671]*kernel[1]+tmp[3672]*kernel[2]+tmp[3770]*kernel[3]+tmp[3771]*kernel[4]+tmp[3772]*kernel[5]+tmp[3870]*kernel[6]+tmp[3871]*kernel[7]+tmp[3872]*kernel[8];
				ans[3772]<=tmp[3671]*kernel[0]+tmp[3672]*kernel[1]+tmp[3673]*kernel[2]+tmp[3771]*kernel[3]+tmp[3772]*kernel[4]+tmp[3773]*kernel[5]+tmp[3871]*kernel[6]+tmp[3872]*kernel[7]+tmp[3873]*kernel[8];
				ans[3773]<=tmp[3672]*kernel[0]+tmp[3673]*kernel[1]+tmp[3674]*kernel[2]+tmp[3772]*kernel[3]+tmp[3773]*kernel[4]+tmp[3774]*kernel[5]+tmp[3872]*kernel[6]+tmp[3873]*kernel[7]+tmp[3874]*kernel[8];
				ans[3774]<=tmp[3673]*kernel[0]+tmp[3674]*kernel[1]+tmp[3675]*kernel[2]+tmp[3773]*kernel[3]+tmp[3774]*kernel[4]+tmp[3775]*kernel[5]+tmp[3873]*kernel[6]+tmp[3874]*kernel[7]+tmp[3875]*kernel[8];
				ans[3775]<=tmp[3674]*kernel[0]+tmp[3675]*kernel[1]+tmp[3676]*kernel[2]+tmp[3774]*kernel[3]+tmp[3775]*kernel[4]+tmp[3776]*kernel[5]+tmp[3874]*kernel[6]+tmp[3875]*kernel[7]+tmp[3876]*kernel[8];
				ans[3776]<=tmp[3675]*kernel[0]+tmp[3676]*kernel[1]+tmp[3677]*kernel[2]+tmp[3775]*kernel[3]+tmp[3776]*kernel[4]+tmp[3777]*kernel[5]+tmp[3875]*kernel[6]+tmp[3876]*kernel[7]+tmp[3877]*kernel[8];
				ans[3777]<=tmp[3676]*kernel[0]+tmp[3677]*kernel[1]+tmp[3678]*kernel[2]+tmp[3776]*kernel[3]+tmp[3777]*kernel[4]+tmp[3778]*kernel[5]+tmp[3876]*kernel[6]+tmp[3877]*kernel[7]+tmp[3878]*kernel[8];
				ans[3778]<=tmp[3677]*kernel[0]+tmp[3678]*kernel[1]+tmp[3679]*kernel[2]+tmp[3777]*kernel[3]+tmp[3778]*kernel[4]+tmp[3779]*kernel[5]+tmp[3877]*kernel[6]+tmp[3878]*kernel[7]+tmp[3879]*kernel[8];
				ans[3779]<=tmp[3678]*kernel[0]+tmp[3679]*kernel[1]+tmp[3680]*kernel[2]+tmp[3778]*kernel[3]+tmp[3779]*kernel[4]+tmp[3780]*kernel[5]+tmp[3878]*kernel[6]+tmp[3879]*kernel[7]+tmp[3880]*kernel[8];
				ans[3780]<=tmp[3679]*kernel[0]+tmp[3680]*kernel[1]+tmp[3681]*kernel[2]+tmp[3779]*kernel[3]+tmp[3780]*kernel[4]+tmp[3781]*kernel[5]+tmp[3879]*kernel[6]+tmp[3880]*kernel[7]+tmp[3881]*kernel[8];
				ans[3781]<=tmp[3680]*kernel[0]+tmp[3681]*kernel[1]+tmp[3682]*kernel[2]+tmp[3780]*kernel[3]+tmp[3781]*kernel[4]+tmp[3782]*kernel[5]+tmp[3880]*kernel[6]+tmp[3881]*kernel[7]+tmp[3882]*kernel[8];
				ans[3782]<=tmp[3681]*kernel[0]+tmp[3682]*kernel[1]+tmp[3683]*kernel[2]+tmp[3781]*kernel[3]+tmp[3782]*kernel[4]+tmp[3783]*kernel[5]+tmp[3881]*kernel[6]+tmp[3882]*kernel[7]+tmp[3883]*kernel[8];
				ans[3783]<=tmp[3682]*kernel[0]+tmp[3683]*kernel[1]+tmp[3684]*kernel[2]+tmp[3782]*kernel[3]+tmp[3783]*kernel[4]+tmp[3784]*kernel[5]+tmp[3882]*kernel[6]+tmp[3883]*kernel[7]+tmp[3884]*kernel[8];
				ans[3784]<=tmp[3683]*kernel[0]+tmp[3684]*kernel[1]+tmp[3685]*kernel[2]+tmp[3783]*kernel[3]+tmp[3784]*kernel[4]+tmp[3785]*kernel[5]+tmp[3883]*kernel[6]+tmp[3884]*kernel[7]+tmp[3885]*kernel[8];
				ans[3785]<=tmp[3684]*kernel[0]+tmp[3685]*kernel[1]+tmp[3686]*kernel[2]+tmp[3784]*kernel[3]+tmp[3785]*kernel[4]+tmp[3786]*kernel[5]+tmp[3884]*kernel[6]+tmp[3885]*kernel[7]+tmp[3886]*kernel[8];
				ans[3786]<=tmp[3685]*kernel[0]+tmp[3686]*kernel[1]+tmp[3687]*kernel[2]+tmp[3785]*kernel[3]+tmp[3786]*kernel[4]+tmp[3787]*kernel[5]+tmp[3885]*kernel[6]+tmp[3886]*kernel[7]+tmp[3887]*kernel[8];
				ans[3787]<=tmp[3686]*kernel[0]+tmp[3687]*kernel[1]+tmp[3688]*kernel[2]+tmp[3786]*kernel[3]+tmp[3787]*kernel[4]+tmp[3788]*kernel[5]+tmp[3886]*kernel[6]+tmp[3887]*kernel[7]+tmp[3888]*kernel[8];
				ans[3788]<=tmp[3687]*kernel[0]+tmp[3688]*kernel[1]+tmp[3689]*kernel[2]+tmp[3787]*kernel[3]+tmp[3788]*kernel[4]+tmp[3789]*kernel[5]+tmp[3887]*kernel[6]+tmp[3888]*kernel[7]+tmp[3889]*kernel[8];
				ans[3789]<=tmp[3688]*kernel[0]+tmp[3689]*kernel[1]+tmp[3690]*kernel[2]+tmp[3788]*kernel[3]+tmp[3789]*kernel[4]+tmp[3790]*kernel[5]+tmp[3888]*kernel[6]+tmp[3889]*kernel[7]+tmp[3890]*kernel[8];
				ans[3790]<=tmp[3689]*kernel[0]+tmp[3690]*kernel[1]+tmp[3691]*kernel[2]+tmp[3789]*kernel[3]+tmp[3790]*kernel[4]+tmp[3791]*kernel[5]+tmp[3889]*kernel[6]+tmp[3890]*kernel[7]+tmp[3891]*kernel[8];
				ans[3791]<=tmp[3690]*kernel[0]+tmp[3691]*kernel[1]+tmp[3692]*kernel[2]+tmp[3790]*kernel[3]+tmp[3791]*kernel[4]+tmp[3792]*kernel[5]+tmp[3890]*kernel[6]+tmp[3891]*kernel[7]+tmp[3892]*kernel[8];
				ans[3792]<=tmp[3691]*kernel[0]+tmp[3692]*kernel[1]+tmp[3693]*kernel[2]+tmp[3791]*kernel[3]+tmp[3792]*kernel[4]+tmp[3793]*kernel[5]+tmp[3891]*kernel[6]+tmp[3892]*kernel[7]+tmp[3893]*kernel[8];
				ans[3793]<=tmp[3692]*kernel[0]+tmp[3693]*kernel[1]+tmp[3694]*kernel[2]+tmp[3792]*kernel[3]+tmp[3793]*kernel[4]+tmp[3794]*kernel[5]+tmp[3892]*kernel[6]+tmp[3893]*kernel[7]+tmp[3894]*kernel[8];
				ans[3794]<=tmp[3693]*kernel[0]+tmp[3694]*kernel[1]+tmp[3695]*kernel[2]+tmp[3793]*kernel[3]+tmp[3794]*kernel[4]+tmp[3795]*kernel[5]+tmp[3893]*kernel[6]+tmp[3894]*kernel[7]+tmp[3895]*kernel[8];
				ans[3795]<=tmp[3694]*kernel[0]+tmp[3695]*kernel[1]+tmp[3696]*kernel[2]+tmp[3794]*kernel[3]+tmp[3795]*kernel[4]+tmp[3796]*kernel[5]+tmp[3894]*kernel[6]+tmp[3895]*kernel[7]+tmp[3896]*kernel[8];
				ans[3796]<=tmp[3695]*kernel[0]+tmp[3696]*kernel[1]+tmp[3697]*kernel[2]+tmp[3795]*kernel[3]+tmp[3796]*kernel[4]+tmp[3797]*kernel[5]+tmp[3895]*kernel[6]+tmp[3896]*kernel[7]+tmp[3897]*kernel[8];
				ans[3797]<=tmp[3696]*kernel[0]+tmp[3697]*kernel[1]+tmp[3698]*kernel[2]+tmp[3796]*kernel[3]+tmp[3797]*kernel[4]+tmp[3798]*kernel[5]+tmp[3896]*kernel[6]+tmp[3897]*kernel[7]+tmp[3898]*kernel[8];
				ans[3798]<=tmp[3697]*kernel[0]+tmp[3698]*kernel[1]+tmp[3699]*kernel[2]+tmp[3797]*kernel[3]+tmp[3798]*kernel[4]+tmp[3799]*kernel[5]+tmp[3897]*kernel[6]+tmp[3898]*kernel[7]+tmp[3899]*kernel[8];
				ans[3799]<=tmp[3698]*kernel[0]+tmp[3699]*kernel[1]+tmp[3798]*kernel[3]+tmp[3799]*kernel[4]+tmp[3898]*kernel[6]+tmp[3899]*kernel[7];
				ans[3800]<=tmp[3700]*kernel[1]+tmp[3701]*kernel[2]+tmp[3800]*kernel[4]+tmp[3801]*kernel[5]+tmp[3900]*kernel[7]+tmp[3901]*kernel[8];
				ans[3801]<=tmp[3700]*kernel[0]+tmp[3701]*kernel[1]+tmp[3702]*kernel[2]+tmp[3800]*kernel[3]+tmp[3801]*kernel[4]+tmp[3802]*kernel[5]+tmp[3900]*kernel[6]+tmp[3901]*kernel[7]+tmp[3902]*kernel[8];
				ans[3802]<=tmp[3701]*kernel[0]+tmp[3702]*kernel[1]+tmp[3703]*kernel[2]+tmp[3801]*kernel[3]+tmp[3802]*kernel[4]+tmp[3803]*kernel[5]+tmp[3901]*kernel[6]+tmp[3902]*kernel[7]+tmp[3903]*kernel[8];
				ans[3803]<=tmp[3702]*kernel[0]+tmp[3703]*kernel[1]+tmp[3704]*kernel[2]+tmp[3802]*kernel[3]+tmp[3803]*kernel[4]+tmp[3804]*kernel[5]+tmp[3902]*kernel[6]+tmp[3903]*kernel[7]+tmp[3904]*kernel[8];
				ans[3804]<=tmp[3703]*kernel[0]+tmp[3704]*kernel[1]+tmp[3705]*kernel[2]+tmp[3803]*kernel[3]+tmp[3804]*kernel[4]+tmp[3805]*kernel[5]+tmp[3903]*kernel[6]+tmp[3904]*kernel[7]+tmp[3905]*kernel[8];
				ans[3805]<=tmp[3704]*kernel[0]+tmp[3705]*kernel[1]+tmp[3706]*kernel[2]+tmp[3804]*kernel[3]+tmp[3805]*kernel[4]+tmp[3806]*kernel[5]+tmp[3904]*kernel[6]+tmp[3905]*kernel[7]+tmp[3906]*kernel[8];
				ans[3806]<=tmp[3705]*kernel[0]+tmp[3706]*kernel[1]+tmp[3707]*kernel[2]+tmp[3805]*kernel[3]+tmp[3806]*kernel[4]+tmp[3807]*kernel[5]+tmp[3905]*kernel[6]+tmp[3906]*kernel[7]+tmp[3907]*kernel[8];
				ans[3807]<=tmp[3706]*kernel[0]+tmp[3707]*kernel[1]+tmp[3708]*kernel[2]+tmp[3806]*kernel[3]+tmp[3807]*kernel[4]+tmp[3808]*kernel[5]+tmp[3906]*kernel[6]+tmp[3907]*kernel[7]+tmp[3908]*kernel[8];
				ans[3808]<=tmp[3707]*kernel[0]+tmp[3708]*kernel[1]+tmp[3709]*kernel[2]+tmp[3807]*kernel[3]+tmp[3808]*kernel[4]+tmp[3809]*kernel[5]+tmp[3907]*kernel[6]+tmp[3908]*kernel[7]+tmp[3909]*kernel[8];
				ans[3809]<=tmp[3708]*kernel[0]+tmp[3709]*kernel[1]+tmp[3710]*kernel[2]+tmp[3808]*kernel[3]+tmp[3809]*kernel[4]+tmp[3810]*kernel[5]+tmp[3908]*kernel[6]+tmp[3909]*kernel[7]+tmp[3910]*kernel[8];
				ans[3810]<=tmp[3709]*kernel[0]+tmp[3710]*kernel[1]+tmp[3711]*kernel[2]+tmp[3809]*kernel[3]+tmp[3810]*kernel[4]+tmp[3811]*kernel[5]+tmp[3909]*kernel[6]+tmp[3910]*kernel[7]+tmp[3911]*kernel[8];
				ans[3811]<=tmp[3710]*kernel[0]+tmp[3711]*kernel[1]+tmp[3712]*kernel[2]+tmp[3810]*kernel[3]+tmp[3811]*kernel[4]+tmp[3812]*kernel[5]+tmp[3910]*kernel[6]+tmp[3911]*kernel[7]+tmp[3912]*kernel[8];
				ans[3812]<=tmp[3711]*kernel[0]+tmp[3712]*kernel[1]+tmp[3713]*kernel[2]+tmp[3811]*kernel[3]+tmp[3812]*kernel[4]+tmp[3813]*kernel[5]+tmp[3911]*kernel[6]+tmp[3912]*kernel[7]+tmp[3913]*kernel[8];
				ans[3813]<=tmp[3712]*kernel[0]+tmp[3713]*kernel[1]+tmp[3714]*kernel[2]+tmp[3812]*kernel[3]+tmp[3813]*kernel[4]+tmp[3814]*kernel[5]+tmp[3912]*kernel[6]+tmp[3913]*kernel[7]+tmp[3914]*kernel[8];
				ans[3814]<=tmp[3713]*kernel[0]+tmp[3714]*kernel[1]+tmp[3715]*kernel[2]+tmp[3813]*kernel[3]+tmp[3814]*kernel[4]+tmp[3815]*kernel[5]+tmp[3913]*kernel[6]+tmp[3914]*kernel[7]+tmp[3915]*kernel[8];
				ans[3815]<=tmp[3714]*kernel[0]+tmp[3715]*kernel[1]+tmp[3716]*kernel[2]+tmp[3814]*kernel[3]+tmp[3815]*kernel[4]+tmp[3816]*kernel[5]+tmp[3914]*kernel[6]+tmp[3915]*kernel[7]+tmp[3916]*kernel[8];
				ans[3816]<=tmp[3715]*kernel[0]+tmp[3716]*kernel[1]+tmp[3717]*kernel[2]+tmp[3815]*kernel[3]+tmp[3816]*kernel[4]+tmp[3817]*kernel[5]+tmp[3915]*kernel[6]+tmp[3916]*kernel[7]+tmp[3917]*kernel[8];
				ans[3817]<=tmp[3716]*kernel[0]+tmp[3717]*kernel[1]+tmp[3718]*kernel[2]+tmp[3816]*kernel[3]+tmp[3817]*kernel[4]+tmp[3818]*kernel[5]+tmp[3916]*kernel[6]+tmp[3917]*kernel[7]+tmp[3918]*kernel[8];
				ans[3818]<=tmp[3717]*kernel[0]+tmp[3718]*kernel[1]+tmp[3719]*kernel[2]+tmp[3817]*kernel[3]+tmp[3818]*kernel[4]+tmp[3819]*kernel[5]+tmp[3917]*kernel[6]+tmp[3918]*kernel[7]+tmp[3919]*kernel[8];
				ans[3819]<=tmp[3718]*kernel[0]+tmp[3719]*kernel[1]+tmp[3720]*kernel[2]+tmp[3818]*kernel[3]+tmp[3819]*kernel[4]+tmp[3820]*kernel[5]+tmp[3918]*kernel[6]+tmp[3919]*kernel[7]+tmp[3920]*kernel[8];
				ans[3820]<=tmp[3719]*kernel[0]+tmp[3720]*kernel[1]+tmp[3721]*kernel[2]+tmp[3819]*kernel[3]+tmp[3820]*kernel[4]+tmp[3821]*kernel[5]+tmp[3919]*kernel[6]+tmp[3920]*kernel[7]+tmp[3921]*kernel[8];
				ans[3821]<=tmp[3720]*kernel[0]+tmp[3721]*kernel[1]+tmp[3722]*kernel[2]+tmp[3820]*kernel[3]+tmp[3821]*kernel[4]+tmp[3822]*kernel[5]+tmp[3920]*kernel[6]+tmp[3921]*kernel[7]+tmp[3922]*kernel[8];
				ans[3822]<=tmp[3721]*kernel[0]+tmp[3722]*kernel[1]+tmp[3723]*kernel[2]+tmp[3821]*kernel[3]+tmp[3822]*kernel[4]+tmp[3823]*kernel[5]+tmp[3921]*kernel[6]+tmp[3922]*kernel[7]+tmp[3923]*kernel[8];
				ans[3823]<=tmp[3722]*kernel[0]+tmp[3723]*kernel[1]+tmp[3724]*kernel[2]+tmp[3822]*kernel[3]+tmp[3823]*kernel[4]+tmp[3824]*kernel[5]+tmp[3922]*kernel[6]+tmp[3923]*kernel[7]+tmp[3924]*kernel[8];
				ans[3824]<=tmp[3723]*kernel[0]+tmp[3724]*kernel[1]+tmp[3725]*kernel[2]+tmp[3823]*kernel[3]+tmp[3824]*kernel[4]+tmp[3825]*kernel[5]+tmp[3923]*kernel[6]+tmp[3924]*kernel[7]+tmp[3925]*kernel[8];
				ans[3825]<=tmp[3724]*kernel[0]+tmp[3725]*kernel[1]+tmp[3726]*kernel[2]+tmp[3824]*kernel[3]+tmp[3825]*kernel[4]+tmp[3826]*kernel[5]+tmp[3924]*kernel[6]+tmp[3925]*kernel[7]+tmp[3926]*kernel[8];
				ans[3826]<=tmp[3725]*kernel[0]+tmp[3726]*kernel[1]+tmp[3727]*kernel[2]+tmp[3825]*kernel[3]+tmp[3826]*kernel[4]+tmp[3827]*kernel[5]+tmp[3925]*kernel[6]+tmp[3926]*kernel[7]+tmp[3927]*kernel[8];
				ans[3827]<=tmp[3726]*kernel[0]+tmp[3727]*kernel[1]+tmp[3728]*kernel[2]+tmp[3826]*kernel[3]+tmp[3827]*kernel[4]+tmp[3828]*kernel[5]+tmp[3926]*kernel[6]+tmp[3927]*kernel[7]+tmp[3928]*kernel[8];
				ans[3828]<=tmp[3727]*kernel[0]+tmp[3728]*kernel[1]+tmp[3729]*kernel[2]+tmp[3827]*kernel[3]+tmp[3828]*kernel[4]+tmp[3829]*kernel[5]+tmp[3927]*kernel[6]+tmp[3928]*kernel[7]+tmp[3929]*kernel[8];
				ans[3829]<=tmp[3728]*kernel[0]+tmp[3729]*kernel[1]+tmp[3730]*kernel[2]+tmp[3828]*kernel[3]+tmp[3829]*kernel[4]+tmp[3830]*kernel[5]+tmp[3928]*kernel[6]+tmp[3929]*kernel[7]+tmp[3930]*kernel[8];
				ans[3830]<=tmp[3729]*kernel[0]+tmp[3730]*kernel[1]+tmp[3731]*kernel[2]+tmp[3829]*kernel[3]+tmp[3830]*kernel[4]+tmp[3831]*kernel[5]+tmp[3929]*kernel[6]+tmp[3930]*kernel[7]+tmp[3931]*kernel[8];
				ans[3831]<=tmp[3730]*kernel[0]+tmp[3731]*kernel[1]+tmp[3732]*kernel[2]+tmp[3830]*kernel[3]+tmp[3831]*kernel[4]+tmp[3832]*kernel[5]+tmp[3930]*kernel[6]+tmp[3931]*kernel[7]+tmp[3932]*kernel[8];
				ans[3832]<=tmp[3731]*kernel[0]+tmp[3732]*kernel[1]+tmp[3733]*kernel[2]+tmp[3831]*kernel[3]+tmp[3832]*kernel[4]+tmp[3833]*kernel[5]+tmp[3931]*kernel[6]+tmp[3932]*kernel[7]+tmp[3933]*kernel[8];
				ans[3833]<=tmp[3732]*kernel[0]+tmp[3733]*kernel[1]+tmp[3734]*kernel[2]+tmp[3832]*kernel[3]+tmp[3833]*kernel[4]+tmp[3834]*kernel[5]+tmp[3932]*kernel[6]+tmp[3933]*kernel[7]+tmp[3934]*kernel[8];
				ans[3834]<=tmp[3733]*kernel[0]+tmp[3734]*kernel[1]+tmp[3735]*kernel[2]+tmp[3833]*kernel[3]+tmp[3834]*kernel[4]+tmp[3835]*kernel[5]+tmp[3933]*kernel[6]+tmp[3934]*kernel[7]+tmp[3935]*kernel[8];
				ans[3835]<=tmp[3734]*kernel[0]+tmp[3735]*kernel[1]+tmp[3736]*kernel[2]+tmp[3834]*kernel[3]+tmp[3835]*kernel[4]+tmp[3836]*kernel[5]+tmp[3934]*kernel[6]+tmp[3935]*kernel[7]+tmp[3936]*kernel[8];
				ans[3836]<=tmp[3735]*kernel[0]+tmp[3736]*kernel[1]+tmp[3737]*kernel[2]+tmp[3835]*kernel[3]+tmp[3836]*kernel[4]+tmp[3837]*kernel[5]+tmp[3935]*kernel[6]+tmp[3936]*kernel[7]+tmp[3937]*kernel[8];
				ans[3837]<=tmp[3736]*kernel[0]+tmp[3737]*kernel[1]+tmp[3738]*kernel[2]+tmp[3836]*kernel[3]+tmp[3837]*kernel[4]+tmp[3838]*kernel[5]+tmp[3936]*kernel[6]+tmp[3937]*kernel[7]+tmp[3938]*kernel[8];
				ans[3838]<=tmp[3737]*kernel[0]+tmp[3738]*kernel[1]+tmp[3739]*kernel[2]+tmp[3837]*kernel[3]+tmp[3838]*kernel[4]+tmp[3839]*kernel[5]+tmp[3937]*kernel[6]+tmp[3938]*kernel[7]+tmp[3939]*kernel[8];
				ans[3839]<=tmp[3738]*kernel[0]+tmp[3739]*kernel[1]+tmp[3740]*kernel[2]+tmp[3838]*kernel[3]+tmp[3839]*kernel[4]+tmp[3840]*kernel[5]+tmp[3938]*kernel[6]+tmp[3939]*kernel[7]+tmp[3940]*kernel[8];
				ans[3840]<=tmp[3739]*kernel[0]+tmp[3740]*kernel[1]+tmp[3741]*kernel[2]+tmp[3839]*kernel[3]+tmp[3840]*kernel[4]+tmp[3841]*kernel[5]+tmp[3939]*kernel[6]+tmp[3940]*kernel[7]+tmp[3941]*kernel[8];
				ans[3841]<=tmp[3740]*kernel[0]+tmp[3741]*kernel[1]+tmp[3742]*kernel[2]+tmp[3840]*kernel[3]+tmp[3841]*kernel[4]+tmp[3842]*kernel[5]+tmp[3940]*kernel[6]+tmp[3941]*kernel[7]+tmp[3942]*kernel[8];
				ans[3842]<=tmp[3741]*kernel[0]+tmp[3742]*kernel[1]+tmp[3743]*kernel[2]+tmp[3841]*kernel[3]+tmp[3842]*kernel[4]+tmp[3843]*kernel[5]+tmp[3941]*kernel[6]+tmp[3942]*kernel[7]+tmp[3943]*kernel[8];
				ans[3843]<=tmp[3742]*kernel[0]+tmp[3743]*kernel[1]+tmp[3744]*kernel[2]+tmp[3842]*kernel[3]+tmp[3843]*kernel[4]+tmp[3844]*kernel[5]+tmp[3942]*kernel[6]+tmp[3943]*kernel[7]+tmp[3944]*kernel[8];
				ans[3844]<=tmp[3743]*kernel[0]+tmp[3744]*kernel[1]+tmp[3745]*kernel[2]+tmp[3843]*kernel[3]+tmp[3844]*kernel[4]+tmp[3845]*kernel[5]+tmp[3943]*kernel[6]+tmp[3944]*kernel[7]+tmp[3945]*kernel[8];
				ans[3845]<=tmp[3744]*kernel[0]+tmp[3745]*kernel[1]+tmp[3746]*kernel[2]+tmp[3844]*kernel[3]+tmp[3845]*kernel[4]+tmp[3846]*kernel[5]+tmp[3944]*kernel[6]+tmp[3945]*kernel[7]+tmp[3946]*kernel[8];
				ans[3846]<=tmp[3745]*kernel[0]+tmp[3746]*kernel[1]+tmp[3747]*kernel[2]+tmp[3845]*kernel[3]+tmp[3846]*kernel[4]+tmp[3847]*kernel[5]+tmp[3945]*kernel[6]+tmp[3946]*kernel[7]+tmp[3947]*kernel[8];
				ans[3847]<=tmp[3746]*kernel[0]+tmp[3747]*kernel[1]+tmp[3748]*kernel[2]+tmp[3846]*kernel[3]+tmp[3847]*kernel[4]+tmp[3848]*kernel[5]+tmp[3946]*kernel[6]+tmp[3947]*kernel[7]+tmp[3948]*kernel[8];
				ans[3848]<=tmp[3747]*kernel[0]+tmp[3748]*kernel[1]+tmp[3749]*kernel[2]+tmp[3847]*kernel[3]+tmp[3848]*kernel[4]+tmp[3849]*kernel[5]+tmp[3947]*kernel[6]+tmp[3948]*kernel[7]+tmp[3949]*kernel[8];
				ans[3849]<=tmp[3748]*kernel[0]+tmp[3749]*kernel[1]+tmp[3750]*kernel[2]+tmp[3848]*kernel[3]+tmp[3849]*kernel[4]+tmp[3850]*kernel[5]+tmp[3948]*kernel[6]+tmp[3949]*kernel[7]+tmp[3950]*kernel[8];
				ans[3850]<=tmp[3749]*kernel[0]+tmp[3750]*kernel[1]+tmp[3751]*kernel[2]+tmp[3849]*kernel[3]+tmp[3850]*kernel[4]+tmp[3851]*kernel[5]+tmp[3949]*kernel[6]+tmp[3950]*kernel[7]+tmp[3951]*kernel[8];
				ans[3851]<=tmp[3750]*kernel[0]+tmp[3751]*kernel[1]+tmp[3752]*kernel[2]+tmp[3850]*kernel[3]+tmp[3851]*kernel[4]+tmp[3852]*kernel[5]+tmp[3950]*kernel[6]+tmp[3951]*kernel[7]+tmp[3952]*kernel[8];
				ans[3852]<=tmp[3751]*kernel[0]+tmp[3752]*kernel[1]+tmp[3753]*kernel[2]+tmp[3851]*kernel[3]+tmp[3852]*kernel[4]+tmp[3853]*kernel[5]+tmp[3951]*kernel[6]+tmp[3952]*kernel[7]+tmp[3953]*kernel[8];
				ans[3853]<=tmp[3752]*kernel[0]+tmp[3753]*kernel[1]+tmp[3754]*kernel[2]+tmp[3852]*kernel[3]+tmp[3853]*kernel[4]+tmp[3854]*kernel[5]+tmp[3952]*kernel[6]+tmp[3953]*kernel[7]+tmp[3954]*kernel[8];
				ans[3854]<=tmp[3753]*kernel[0]+tmp[3754]*kernel[1]+tmp[3755]*kernel[2]+tmp[3853]*kernel[3]+tmp[3854]*kernel[4]+tmp[3855]*kernel[5]+tmp[3953]*kernel[6]+tmp[3954]*kernel[7]+tmp[3955]*kernel[8];
				ans[3855]<=tmp[3754]*kernel[0]+tmp[3755]*kernel[1]+tmp[3756]*kernel[2]+tmp[3854]*kernel[3]+tmp[3855]*kernel[4]+tmp[3856]*kernel[5]+tmp[3954]*kernel[6]+tmp[3955]*kernel[7]+tmp[3956]*kernel[8];
				ans[3856]<=tmp[3755]*kernel[0]+tmp[3756]*kernel[1]+tmp[3757]*kernel[2]+tmp[3855]*kernel[3]+tmp[3856]*kernel[4]+tmp[3857]*kernel[5]+tmp[3955]*kernel[6]+tmp[3956]*kernel[7]+tmp[3957]*kernel[8];
				ans[3857]<=tmp[3756]*kernel[0]+tmp[3757]*kernel[1]+tmp[3758]*kernel[2]+tmp[3856]*kernel[3]+tmp[3857]*kernel[4]+tmp[3858]*kernel[5]+tmp[3956]*kernel[6]+tmp[3957]*kernel[7]+tmp[3958]*kernel[8];
				ans[3858]<=tmp[3757]*kernel[0]+tmp[3758]*kernel[1]+tmp[3759]*kernel[2]+tmp[3857]*kernel[3]+tmp[3858]*kernel[4]+tmp[3859]*kernel[5]+tmp[3957]*kernel[6]+tmp[3958]*kernel[7]+tmp[3959]*kernel[8];
				ans[3859]<=tmp[3758]*kernel[0]+tmp[3759]*kernel[1]+tmp[3760]*kernel[2]+tmp[3858]*kernel[3]+tmp[3859]*kernel[4]+tmp[3860]*kernel[5]+tmp[3958]*kernel[6]+tmp[3959]*kernel[7]+tmp[3960]*kernel[8];
				ans[3860]<=tmp[3759]*kernel[0]+tmp[3760]*kernel[1]+tmp[3761]*kernel[2]+tmp[3859]*kernel[3]+tmp[3860]*kernel[4]+tmp[3861]*kernel[5]+tmp[3959]*kernel[6]+tmp[3960]*kernel[7]+tmp[3961]*kernel[8];
				ans[3861]<=tmp[3760]*kernel[0]+tmp[3761]*kernel[1]+tmp[3762]*kernel[2]+tmp[3860]*kernel[3]+tmp[3861]*kernel[4]+tmp[3862]*kernel[5]+tmp[3960]*kernel[6]+tmp[3961]*kernel[7]+tmp[3962]*kernel[8];
				ans[3862]<=tmp[3761]*kernel[0]+tmp[3762]*kernel[1]+tmp[3763]*kernel[2]+tmp[3861]*kernel[3]+tmp[3862]*kernel[4]+tmp[3863]*kernel[5]+tmp[3961]*kernel[6]+tmp[3962]*kernel[7]+tmp[3963]*kernel[8];
				ans[3863]<=tmp[3762]*kernel[0]+tmp[3763]*kernel[1]+tmp[3764]*kernel[2]+tmp[3862]*kernel[3]+tmp[3863]*kernel[4]+tmp[3864]*kernel[5]+tmp[3962]*kernel[6]+tmp[3963]*kernel[7]+tmp[3964]*kernel[8];
				ans[3864]<=tmp[3763]*kernel[0]+tmp[3764]*kernel[1]+tmp[3765]*kernel[2]+tmp[3863]*kernel[3]+tmp[3864]*kernel[4]+tmp[3865]*kernel[5]+tmp[3963]*kernel[6]+tmp[3964]*kernel[7]+tmp[3965]*kernel[8];
				ans[3865]<=tmp[3764]*kernel[0]+tmp[3765]*kernel[1]+tmp[3766]*kernel[2]+tmp[3864]*kernel[3]+tmp[3865]*kernel[4]+tmp[3866]*kernel[5]+tmp[3964]*kernel[6]+tmp[3965]*kernel[7]+tmp[3966]*kernel[8];
				ans[3866]<=tmp[3765]*kernel[0]+tmp[3766]*kernel[1]+tmp[3767]*kernel[2]+tmp[3865]*kernel[3]+tmp[3866]*kernel[4]+tmp[3867]*kernel[5]+tmp[3965]*kernel[6]+tmp[3966]*kernel[7]+tmp[3967]*kernel[8];
				ans[3867]<=tmp[3766]*kernel[0]+tmp[3767]*kernel[1]+tmp[3768]*kernel[2]+tmp[3866]*kernel[3]+tmp[3867]*kernel[4]+tmp[3868]*kernel[5]+tmp[3966]*kernel[6]+tmp[3967]*kernel[7]+tmp[3968]*kernel[8];
				ans[3868]<=tmp[3767]*kernel[0]+tmp[3768]*kernel[1]+tmp[3769]*kernel[2]+tmp[3867]*kernel[3]+tmp[3868]*kernel[4]+tmp[3869]*kernel[5]+tmp[3967]*kernel[6]+tmp[3968]*kernel[7]+tmp[3969]*kernel[8];
				ans[3869]<=tmp[3768]*kernel[0]+tmp[3769]*kernel[1]+tmp[3770]*kernel[2]+tmp[3868]*kernel[3]+tmp[3869]*kernel[4]+tmp[3870]*kernel[5]+tmp[3968]*kernel[6]+tmp[3969]*kernel[7]+tmp[3970]*kernel[8];
				ans[3870]<=tmp[3769]*kernel[0]+tmp[3770]*kernel[1]+tmp[3771]*kernel[2]+tmp[3869]*kernel[3]+tmp[3870]*kernel[4]+tmp[3871]*kernel[5]+tmp[3969]*kernel[6]+tmp[3970]*kernel[7]+tmp[3971]*kernel[8];
				ans[3871]<=tmp[3770]*kernel[0]+tmp[3771]*kernel[1]+tmp[3772]*kernel[2]+tmp[3870]*kernel[3]+tmp[3871]*kernel[4]+tmp[3872]*kernel[5]+tmp[3970]*kernel[6]+tmp[3971]*kernel[7]+tmp[3972]*kernel[8];
				ans[3872]<=tmp[3771]*kernel[0]+tmp[3772]*kernel[1]+tmp[3773]*kernel[2]+tmp[3871]*kernel[3]+tmp[3872]*kernel[4]+tmp[3873]*kernel[5]+tmp[3971]*kernel[6]+tmp[3972]*kernel[7]+tmp[3973]*kernel[8];
				ans[3873]<=tmp[3772]*kernel[0]+tmp[3773]*kernel[1]+tmp[3774]*kernel[2]+tmp[3872]*kernel[3]+tmp[3873]*kernel[4]+tmp[3874]*kernel[5]+tmp[3972]*kernel[6]+tmp[3973]*kernel[7]+tmp[3974]*kernel[8];
				ans[3874]<=tmp[3773]*kernel[0]+tmp[3774]*kernel[1]+tmp[3775]*kernel[2]+tmp[3873]*kernel[3]+tmp[3874]*kernel[4]+tmp[3875]*kernel[5]+tmp[3973]*kernel[6]+tmp[3974]*kernel[7]+tmp[3975]*kernel[8];
				ans[3875]<=tmp[3774]*kernel[0]+tmp[3775]*kernel[1]+tmp[3776]*kernel[2]+tmp[3874]*kernel[3]+tmp[3875]*kernel[4]+tmp[3876]*kernel[5]+tmp[3974]*kernel[6]+tmp[3975]*kernel[7]+tmp[3976]*kernel[8];
				ans[3876]<=tmp[3775]*kernel[0]+tmp[3776]*kernel[1]+tmp[3777]*kernel[2]+tmp[3875]*kernel[3]+tmp[3876]*kernel[4]+tmp[3877]*kernel[5]+tmp[3975]*kernel[6]+tmp[3976]*kernel[7]+tmp[3977]*kernel[8];
				ans[3877]<=tmp[3776]*kernel[0]+tmp[3777]*kernel[1]+tmp[3778]*kernel[2]+tmp[3876]*kernel[3]+tmp[3877]*kernel[4]+tmp[3878]*kernel[5]+tmp[3976]*kernel[6]+tmp[3977]*kernel[7]+tmp[3978]*kernel[8];
				ans[3878]<=tmp[3777]*kernel[0]+tmp[3778]*kernel[1]+tmp[3779]*kernel[2]+tmp[3877]*kernel[3]+tmp[3878]*kernel[4]+tmp[3879]*kernel[5]+tmp[3977]*kernel[6]+tmp[3978]*kernel[7]+tmp[3979]*kernel[8];
				ans[3879]<=tmp[3778]*kernel[0]+tmp[3779]*kernel[1]+tmp[3780]*kernel[2]+tmp[3878]*kernel[3]+tmp[3879]*kernel[4]+tmp[3880]*kernel[5]+tmp[3978]*kernel[6]+tmp[3979]*kernel[7]+tmp[3980]*kernel[8];
				ans[3880]<=tmp[3779]*kernel[0]+tmp[3780]*kernel[1]+tmp[3781]*kernel[2]+tmp[3879]*kernel[3]+tmp[3880]*kernel[4]+tmp[3881]*kernel[5]+tmp[3979]*kernel[6]+tmp[3980]*kernel[7]+tmp[3981]*kernel[8];
				ans[3881]<=tmp[3780]*kernel[0]+tmp[3781]*kernel[1]+tmp[3782]*kernel[2]+tmp[3880]*kernel[3]+tmp[3881]*kernel[4]+tmp[3882]*kernel[5]+tmp[3980]*kernel[6]+tmp[3981]*kernel[7]+tmp[3982]*kernel[8];
				ans[3882]<=tmp[3781]*kernel[0]+tmp[3782]*kernel[1]+tmp[3783]*kernel[2]+tmp[3881]*kernel[3]+tmp[3882]*kernel[4]+tmp[3883]*kernel[5]+tmp[3981]*kernel[6]+tmp[3982]*kernel[7]+tmp[3983]*kernel[8];
				ans[3883]<=tmp[3782]*kernel[0]+tmp[3783]*kernel[1]+tmp[3784]*kernel[2]+tmp[3882]*kernel[3]+tmp[3883]*kernel[4]+tmp[3884]*kernel[5]+tmp[3982]*kernel[6]+tmp[3983]*kernel[7]+tmp[3984]*kernel[8];
				ans[3884]<=tmp[3783]*kernel[0]+tmp[3784]*kernel[1]+tmp[3785]*kernel[2]+tmp[3883]*kernel[3]+tmp[3884]*kernel[4]+tmp[3885]*kernel[5]+tmp[3983]*kernel[6]+tmp[3984]*kernel[7]+tmp[3985]*kernel[8];
				ans[3885]<=tmp[3784]*kernel[0]+tmp[3785]*kernel[1]+tmp[3786]*kernel[2]+tmp[3884]*kernel[3]+tmp[3885]*kernel[4]+tmp[3886]*kernel[5]+tmp[3984]*kernel[6]+tmp[3985]*kernel[7]+tmp[3986]*kernel[8];
				ans[3886]<=tmp[3785]*kernel[0]+tmp[3786]*kernel[1]+tmp[3787]*kernel[2]+tmp[3885]*kernel[3]+tmp[3886]*kernel[4]+tmp[3887]*kernel[5]+tmp[3985]*kernel[6]+tmp[3986]*kernel[7]+tmp[3987]*kernel[8];
				ans[3887]<=tmp[3786]*kernel[0]+tmp[3787]*kernel[1]+tmp[3788]*kernel[2]+tmp[3886]*kernel[3]+tmp[3887]*kernel[4]+tmp[3888]*kernel[5]+tmp[3986]*kernel[6]+tmp[3987]*kernel[7]+tmp[3988]*kernel[8];
				ans[3888]<=tmp[3787]*kernel[0]+tmp[3788]*kernel[1]+tmp[3789]*kernel[2]+tmp[3887]*kernel[3]+tmp[3888]*kernel[4]+tmp[3889]*kernel[5]+tmp[3987]*kernel[6]+tmp[3988]*kernel[7]+tmp[3989]*kernel[8];
				ans[3889]<=tmp[3788]*kernel[0]+tmp[3789]*kernel[1]+tmp[3790]*kernel[2]+tmp[3888]*kernel[3]+tmp[3889]*kernel[4]+tmp[3890]*kernel[5]+tmp[3988]*kernel[6]+tmp[3989]*kernel[7]+tmp[3990]*kernel[8];
				ans[3890]<=tmp[3789]*kernel[0]+tmp[3790]*kernel[1]+tmp[3791]*kernel[2]+tmp[3889]*kernel[3]+tmp[3890]*kernel[4]+tmp[3891]*kernel[5]+tmp[3989]*kernel[6]+tmp[3990]*kernel[7]+tmp[3991]*kernel[8];
				ans[3891]<=tmp[3790]*kernel[0]+tmp[3791]*kernel[1]+tmp[3792]*kernel[2]+tmp[3890]*kernel[3]+tmp[3891]*kernel[4]+tmp[3892]*kernel[5]+tmp[3990]*kernel[6]+tmp[3991]*kernel[7]+tmp[3992]*kernel[8];
				ans[3892]<=tmp[3791]*kernel[0]+tmp[3792]*kernel[1]+tmp[3793]*kernel[2]+tmp[3891]*kernel[3]+tmp[3892]*kernel[4]+tmp[3893]*kernel[5]+tmp[3991]*kernel[6]+tmp[3992]*kernel[7]+tmp[3993]*kernel[8];
				ans[3893]<=tmp[3792]*kernel[0]+tmp[3793]*kernel[1]+tmp[3794]*kernel[2]+tmp[3892]*kernel[3]+tmp[3893]*kernel[4]+tmp[3894]*kernel[5]+tmp[3992]*kernel[6]+tmp[3993]*kernel[7]+tmp[3994]*kernel[8];
				ans[3894]<=tmp[3793]*kernel[0]+tmp[3794]*kernel[1]+tmp[3795]*kernel[2]+tmp[3893]*kernel[3]+tmp[3894]*kernel[4]+tmp[3895]*kernel[5]+tmp[3993]*kernel[6]+tmp[3994]*kernel[7]+tmp[3995]*kernel[8];
				ans[3895]<=tmp[3794]*kernel[0]+tmp[3795]*kernel[1]+tmp[3796]*kernel[2]+tmp[3894]*kernel[3]+tmp[3895]*kernel[4]+tmp[3896]*kernel[5]+tmp[3994]*kernel[6]+tmp[3995]*kernel[7]+tmp[3996]*kernel[8];
				ans[3896]<=tmp[3795]*kernel[0]+tmp[3796]*kernel[1]+tmp[3797]*kernel[2]+tmp[3895]*kernel[3]+tmp[3896]*kernel[4]+tmp[3897]*kernel[5]+tmp[3995]*kernel[6]+tmp[3996]*kernel[7]+tmp[3997]*kernel[8];
				ans[3897]<=tmp[3796]*kernel[0]+tmp[3797]*kernel[1]+tmp[3798]*kernel[2]+tmp[3896]*kernel[3]+tmp[3897]*kernel[4]+tmp[3898]*kernel[5]+tmp[3996]*kernel[6]+tmp[3997]*kernel[7]+tmp[3998]*kernel[8];
				ans[3898]<=tmp[3797]*kernel[0]+tmp[3798]*kernel[1]+tmp[3799]*kernel[2]+tmp[3897]*kernel[3]+tmp[3898]*kernel[4]+tmp[3899]*kernel[5]+tmp[3997]*kernel[6]+tmp[3998]*kernel[7]+tmp[3999]*kernel[8];
				ans[3899]<=tmp[3798]*kernel[0]+tmp[3799]*kernel[1]+tmp[3898]*kernel[3]+tmp[3899]*kernel[4]+tmp[3998]*kernel[6]+tmp[3999]*kernel[7];
				ans[3900]<=tmp[3800]*kernel[1]+tmp[3801]*kernel[2]+tmp[3900]*kernel[4]+tmp[3901]*kernel[5]+tmp[4000]*kernel[7]+tmp[4001]*kernel[8];
				ans[3901]<=tmp[3800]*kernel[0]+tmp[3801]*kernel[1]+tmp[3802]*kernel[2]+tmp[3900]*kernel[3]+tmp[3901]*kernel[4]+tmp[3902]*kernel[5]+tmp[4000]*kernel[6]+tmp[4001]*kernel[7]+tmp[4002]*kernel[8];
				ans[3902]<=tmp[3801]*kernel[0]+tmp[3802]*kernel[1]+tmp[3803]*kernel[2]+tmp[3901]*kernel[3]+tmp[3902]*kernel[4]+tmp[3903]*kernel[5]+tmp[4001]*kernel[6]+tmp[4002]*kernel[7]+tmp[4003]*kernel[8];
				ans[3903]<=tmp[3802]*kernel[0]+tmp[3803]*kernel[1]+tmp[3804]*kernel[2]+tmp[3902]*kernel[3]+tmp[3903]*kernel[4]+tmp[3904]*kernel[5]+tmp[4002]*kernel[6]+tmp[4003]*kernel[7]+tmp[4004]*kernel[8];
				ans[3904]<=tmp[3803]*kernel[0]+tmp[3804]*kernel[1]+tmp[3805]*kernel[2]+tmp[3903]*kernel[3]+tmp[3904]*kernel[4]+tmp[3905]*kernel[5]+tmp[4003]*kernel[6]+tmp[4004]*kernel[7]+tmp[4005]*kernel[8];
				ans[3905]<=tmp[3804]*kernel[0]+tmp[3805]*kernel[1]+tmp[3806]*kernel[2]+tmp[3904]*kernel[3]+tmp[3905]*kernel[4]+tmp[3906]*kernel[5]+tmp[4004]*kernel[6]+tmp[4005]*kernel[7]+tmp[4006]*kernel[8];
				ans[3906]<=tmp[3805]*kernel[0]+tmp[3806]*kernel[1]+tmp[3807]*kernel[2]+tmp[3905]*kernel[3]+tmp[3906]*kernel[4]+tmp[3907]*kernel[5]+tmp[4005]*kernel[6]+tmp[4006]*kernel[7]+tmp[4007]*kernel[8];
				ans[3907]<=tmp[3806]*kernel[0]+tmp[3807]*kernel[1]+tmp[3808]*kernel[2]+tmp[3906]*kernel[3]+tmp[3907]*kernel[4]+tmp[3908]*kernel[5]+tmp[4006]*kernel[6]+tmp[4007]*kernel[7]+tmp[4008]*kernel[8];
				ans[3908]<=tmp[3807]*kernel[0]+tmp[3808]*kernel[1]+tmp[3809]*kernel[2]+tmp[3907]*kernel[3]+tmp[3908]*kernel[4]+tmp[3909]*kernel[5]+tmp[4007]*kernel[6]+tmp[4008]*kernel[7]+tmp[4009]*kernel[8];
				ans[3909]<=tmp[3808]*kernel[0]+tmp[3809]*kernel[1]+tmp[3810]*kernel[2]+tmp[3908]*kernel[3]+tmp[3909]*kernel[4]+tmp[3910]*kernel[5]+tmp[4008]*kernel[6]+tmp[4009]*kernel[7]+tmp[4010]*kernel[8];
				ans[3910]<=tmp[3809]*kernel[0]+tmp[3810]*kernel[1]+tmp[3811]*kernel[2]+tmp[3909]*kernel[3]+tmp[3910]*kernel[4]+tmp[3911]*kernel[5]+tmp[4009]*kernel[6]+tmp[4010]*kernel[7]+tmp[4011]*kernel[8];
				ans[3911]<=tmp[3810]*kernel[0]+tmp[3811]*kernel[1]+tmp[3812]*kernel[2]+tmp[3910]*kernel[3]+tmp[3911]*kernel[4]+tmp[3912]*kernel[5]+tmp[4010]*kernel[6]+tmp[4011]*kernel[7]+tmp[4012]*kernel[8];
				ans[3912]<=tmp[3811]*kernel[0]+tmp[3812]*kernel[1]+tmp[3813]*kernel[2]+tmp[3911]*kernel[3]+tmp[3912]*kernel[4]+tmp[3913]*kernel[5]+tmp[4011]*kernel[6]+tmp[4012]*kernel[7]+tmp[4013]*kernel[8];
				ans[3913]<=tmp[3812]*kernel[0]+tmp[3813]*kernel[1]+tmp[3814]*kernel[2]+tmp[3912]*kernel[3]+tmp[3913]*kernel[4]+tmp[3914]*kernel[5]+tmp[4012]*kernel[6]+tmp[4013]*kernel[7]+tmp[4014]*kernel[8];
				ans[3914]<=tmp[3813]*kernel[0]+tmp[3814]*kernel[1]+tmp[3815]*kernel[2]+tmp[3913]*kernel[3]+tmp[3914]*kernel[4]+tmp[3915]*kernel[5]+tmp[4013]*kernel[6]+tmp[4014]*kernel[7]+tmp[4015]*kernel[8];
				ans[3915]<=tmp[3814]*kernel[0]+tmp[3815]*kernel[1]+tmp[3816]*kernel[2]+tmp[3914]*kernel[3]+tmp[3915]*kernel[4]+tmp[3916]*kernel[5]+tmp[4014]*kernel[6]+tmp[4015]*kernel[7]+tmp[4016]*kernel[8];
				ans[3916]<=tmp[3815]*kernel[0]+tmp[3816]*kernel[1]+tmp[3817]*kernel[2]+tmp[3915]*kernel[3]+tmp[3916]*kernel[4]+tmp[3917]*kernel[5]+tmp[4015]*kernel[6]+tmp[4016]*kernel[7]+tmp[4017]*kernel[8];
				ans[3917]<=tmp[3816]*kernel[0]+tmp[3817]*kernel[1]+tmp[3818]*kernel[2]+tmp[3916]*kernel[3]+tmp[3917]*kernel[4]+tmp[3918]*kernel[5]+tmp[4016]*kernel[6]+tmp[4017]*kernel[7]+tmp[4018]*kernel[8];
				ans[3918]<=tmp[3817]*kernel[0]+tmp[3818]*kernel[1]+tmp[3819]*kernel[2]+tmp[3917]*kernel[3]+tmp[3918]*kernel[4]+tmp[3919]*kernel[5]+tmp[4017]*kernel[6]+tmp[4018]*kernel[7]+tmp[4019]*kernel[8];
				ans[3919]<=tmp[3818]*kernel[0]+tmp[3819]*kernel[1]+tmp[3820]*kernel[2]+tmp[3918]*kernel[3]+tmp[3919]*kernel[4]+tmp[3920]*kernel[5]+tmp[4018]*kernel[6]+tmp[4019]*kernel[7]+tmp[4020]*kernel[8];
				ans[3920]<=tmp[3819]*kernel[0]+tmp[3820]*kernel[1]+tmp[3821]*kernel[2]+tmp[3919]*kernel[3]+tmp[3920]*kernel[4]+tmp[3921]*kernel[5]+tmp[4019]*kernel[6]+tmp[4020]*kernel[7]+tmp[4021]*kernel[8];
				ans[3921]<=tmp[3820]*kernel[0]+tmp[3821]*kernel[1]+tmp[3822]*kernel[2]+tmp[3920]*kernel[3]+tmp[3921]*kernel[4]+tmp[3922]*kernel[5]+tmp[4020]*kernel[6]+tmp[4021]*kernel[7]+tmp[4022]*kernel[8];
				ans[3922]<=tmp[3821]*kernel[0]+tmp[3822]*kernel[1]+tmp[3823]*kernel[2]+tmp[3921]*kernel[3]+tmp[3922]*kernel[4]+tmp[3923]*kernel[5]+tmp[4021]*kernel[6]+tmp[4022]*kernel[7]+tmp[4023]*kernel[8];
				ans[3923]<=tmp[3822]*kernel[0]+tmp[3823]*kernel[1]+tmp[3824]*kernel[2]+tmp[3922]*kernel[3]+tmp[3923]*kernel[4]+tmp[3924]*kernel[5]+tmp[4022]*kernel[6]+tmp[4023]*kernel[7]+tmp[4024]*kernel[8];
				ans[3924]<=tmp[3823]*kernel[0]+tmp[3824]*kernel[1]+tmp[3825]*kernel[2]+tmp[3923]*kernel[3]+tmp[3924]*kernel[4]+tmp[3925]*kernel[5]+tmp[4023]*kernel[6]+tmp[4024]*kernel[7]+tmp[4025]*kernel[8];
				ans[3925]<=tmp[3824]*kernel[0]+tmp[3825]*kernel[1]+tmp[3826]*kernel[2]+tmp[3924]*kernel[3]+tmp[3925]*kernel[4]+tmp[3926]*kernel[5]+tmp[4024]*kernel[6]+tmp[4025]*kernel[7]+tmp[4026]*kernel[8];
				ans[3926]<=tmp[3825]*kernel[0]+tmp[3826]*kernel[1]+tmp[3827]*kernel[2]+tmp[3925]*kernel[3]+tmp[3926]*kernel[4]+tmp[3927]*kernel[5]+tmp[4025]*kernel[6]+tmp[4026]*kernel[7]+tmp[4027]*kernel[8];
				ans[3927]<=tmp[3826]*kernel[0]+tmp[3827]*kernel[1]+tmp[3828]*kernel[2]+tmp[3926]*kernel[3]+tmp[3927]*kernel[4]+tmp[3928]*kernel[5]+tmp[4026]*kernel[6]+tmp[4027]*kernel[7]+tmp[4028]*kernel[8];
				ans[3928]<=tmp[3827]*kernel[0]+tmp[3828]*kernel[1]+tmp[3829]*kernel[2]+tmp[3927]*kernel[3]+tmp[3928]*kernel[4]+tmp[3929]*kernel[5]+tmp[4027]*kernel[6]+tmp[4028]*kernel[7]+tmp[4029]*kernel[8];
				ans[3929]<=tmp[3828]*kernel[0]+tmp[3829]*kernel[1]+tmp[3830]*kernel[2]+tmp[3928]*kernel[3]+tmp[3929]*kernel[4]+tmp[3930]*kernel[5]+tmp[4028]*kernel[6]+tmp[4029]*kernel[7]+tmp[4030]*kernel[8];
				ans[3930]<=tmp[3829]*kernel[0]+tmp[3830]*kernel[1]+tmp[3831]*kernel[2]+tmp[3929]*kernel[3]+tmp[3930]*kernel[4]+tmp[3931]*kernel[5]+tmp[4029]*kernel[6]+tmp[4030]*kernel[7]+tmp[4031]*kernel[8];
				ans[3931]<=tmp[3830]*kernel[0]+tmp[3831]*kernel[1]+tmp[3832]*kernel[2]+tmp[3930]*kernel[3]+tmp[3931]*kernel[4]+tmp[3932]*kernel[5]+tmp[4030]*kernel[6]+tmp[4031]*kernel[7]+tmp[4032]*kernel[8];
				ans[3932]<=tmp[3831]*kernel[0]+tmp[3832]*kernel[1]+tmp[3833]*kernel[2]+tmp[3931]*kernel[3]+tmp[3932]*kernel[4]+tmp[3933]*kernel[5]+tmp[4031]*kernel[6]+tmp[4032]*kernel[7]+tmp[4033]*kernel[8];
				ans[3933]<=tmp[3832]*kernel[0]+tmp[3833]*kernel[1]+tmp[3834]*kernel[2]+tmp[3932]*kernel[3]+tmp[3933]*kernel[4]+tmp[3934]*kernel[5]+tmp[4032]*kernel[6]+tmp[4033]*kernel[7]+tmp[4034]*kernel[8];
				ans[3934]<=tmp[3833]*kernel[0]+tmp[3834]*kernel[1]+tmp[3835]*kernel[2]+tmp[3933]*kernel[3]+tmp[3934]*kernel[4]+tmp[3935]*kernel[5]+tmp[4033]*kernel[6]+tmp[4034]*kernel[7]+tmp[4035]*kernel[8];
				ans[3935]<=tmp[3834]*kernel[0]+tmp[3835]*kernel[1]+tmp[3836]*kernel[2]+tmp[3934]*kernel[3]+tmp[3935]*kernel[4]+tmp[3936]*kernel[5]+tmp[4034]*kernel[6]+tmp[4035]*kernel[7]+tmp[4036]*kernel[8];
				ans[3936]<=tmp[3835]*kernel[0]+tmp[3836]*kernel[1]+tmp[3837]*kernel[2]+tmp[3935]*kernel[3]+tmp[3936]*kernel[4]+tmp[3937]*kernel[5]+tmp[4035]*kernel[6]+tmp[4036]*kernel[7]+tmp[4037]*kernel[8];
				ans[3937]<=tmp[3836]*kernel[0]+tmp[3837]*kernel[1]+tmp[3838]*kernel[2]+tmp[3936]*kernel[3]+tmp[3937]*kernel[4]+tmp[3938]*kernel[5]+tmp[4036]*kernel[6]+tmp[4037]*kernel[7]+tmp[4038]*kernel[8];
				ans[3938]<=tmp[3837]*kernel[0]+tmp[3838]*kernel[1]+tmp[3839]*kernel[2]+tmp[3937]*kernel[3]+tmp[3938]*kernel[4]+tmp[3939]*kernel[5]+tmp[4037]*kernel[6]+tmp[4038]*kernel[7]+tmp[4039]*kernel[8];
				ans[3939]<=tmp[3838]*kernel[0]+tmp[3839]*kernel[1]+tmp[3840]*kernel[2]+tmp[3938]*kernel[3]+tmp[3939]*kernel[4]+tmp[3940]*kernel[5]+tmp[4038]*kernel[6]+tmp[4039]*kernel[7]+tmp[4040]*kernel[8];
				ans[3940]<=tmp[3839]*kernel[0]+tmp[3840]*kernel[1]+tmp[3841]*kernel[2]+tmp[3939]*kernel[3]+tmp[3940]*kernel[4]+tmp[3941]*kernel[5]+tmp[4039]*kernel[6]+tmp[4040]*kernel[7]+tmp[4041]*kernel[8];
				ans[3941]<=tmp[3840]*kernel[0]+tmp[3841]*kernel[1]+tmp[3842]*kernel[2]+tmp[3940]*kernel[3]+tmp[3941]*kernel[4]+tmp[3942]*kernel[5]+tmp[4040]*kernel[6]+tmp[4041]*kernel[7]+tmp[4042]*kernel[8];
				ans[3942]<=tmp[3841]*kernel[0]+tmp[3842]*kernel[1]+tmp[3843]*kernel[2]+tmp[3941]*kernel[3]+tmp[3942]*kernel[4]+tmp[3943]*kernel[5]+tmp[4041]*kernel[6]+tmp[4042]*kernel[7]+tmp[4043]*kernel[8];
				ans[3943]<=tmp[3842]*kernel[0]+tmp[3843]*kernel[1]+tmp[3844]*kernel[2]+tmp[3942]*kernel[3]+tmp[3943]*kernel[4]+tmp[3944]*kernel[5]+tmp[4042]*kernel[6]+tmp[4043]*kernel[7]+tmp[4044]*kernel[8];
				ans[3944]<=tmp[3843]*kernel[0]+tmp[3844]*kernel[1]+tmp[3845]*kernel[2]+tmp[3943]*kernel[3]+tmp[3944]*kernel[4]+tmp[3945]*kernel[5]+tmp[4043]*kernel[6]+tmp[4044]*kernel[7]+tmp[4045]*kernel[8];
				ans[3945]<=tmp[3844]*kernel[0]+tmp[3845]*kernel[1]+tmp[3846]*kernel[2]+tmp[3944]*kernel[3]+tmp[3945]*kernel[4]+tmp[3946]*kernel[5]+tmp[4044]*kernel[6]+tmp[4045]*kernel[7]+tmp[4046]*kernel[8];
				ans[3946]<=tmp[3845]*kernel[0]+tmp[3846]*kernel[1]+tmp[3847]*kernel[2]+tmp[3945]*kernel[3]+tmp[3946]*kernel[4]+tmp[3947]*kernel[5]+tmp[4045]*kernel[6]+tmp[4046]*kernel[7]+tmp[4047]*kernel[8];
				ans[3947]<=tmp[3846]*kernel[0]+tmp[3847]*kernel[1]+tmp[3848]*kernel[2]+tmp[3946]*kernel[3]+tmp[3947]*kernel[4]+tmp[3948]*kernel[5]+tmp[4046]*kernel[6]+tmp[4047]*kernel[7]+tmp[4048]*kernel[8];
				ans[3948]<=tmp[3847]*kernel[0]+tmp[3848]*kernel[1]+tmp[3849]*kernel[2]+tmp[3947]*kernel[3]+tmp[3948]*kernel[4]+tmp[3949]*kernel[5]+tmp[4047]*kernel[6]+tmp[4048]*kernel[7]+tmp[4049]*kernel[8];
				ans[3949]<=tmp[3848]*kernel[0]+tmp[3849]*kernel[1]+tmp[3850]*kernel[2]+tmp[3948]*kernel[3]+tmp[3949]*kernel[4]+tmp[3950]*kernel[5]+tmp[4048]*kernel[6]+tmp[4049]*kernel[7]+tmp[4050]*kernel[8];
				ans[3950]<=tmp[3849]*kernel[0]+tmp[3850]*kernel[1]+tmp[3851]*kernel[2]+tmp[3949]*kernel[3]+tmp[3950]*kernel[4]+tmp[3951]*kernel[5]+tmp[4049]*kernel[6]+tmp[4050]*kernel[7]+tmp[4051]*kernel[8];
				ans[3951]<=tmp[3850]*kernel[0]+tmp[3851]*kernel[1]+tmp[3852]*kernel[2]+tmp[3950]*kernel[3]+tmp[3951]*kernel[4]+tmp[3952]*kernel[5]+tmp[4050]*kernel[6]+tmp[4051]*kernel[7]+tmp[4052]*kernel[8];
				ans[3952]<=tmp[3851]*kernel[0]+tmp[3852]*kernel[1]+tmp[3853]*kernel[2]+tmp[3951]*kernel[3]+tmp[3952]*kernel[4]+tmp[3953]*kernel[5]+tmp[4051]*kernel[6]+tmp[4052]*kernel[7]+tmp[4053]*kernel[8];
				ans[3953]<=tmp[3852]*kernel[0]+tmp[3853]*kernel[1]+tmp[3854]*kernel[2]+tmp[3952]*kernel[3]+tmp[3953]*kernel[4]+tmp[3954]*kernel[5]+tmp[4052]*kernel[6]+tmp[4053]*kernel[7]+tmp[4054]*kernel[8];
				ans[3954]<=tmp[3853]*kernel[0]+tmp[3854]*kernel[1]+tmp[3855]*kernel[2]+tmp[3953]*kernel[3]+tmp[3954]*kernel[4]+tmp[3955]*kernel[5]+tmp[4053]*kernel[6]+tmp[4054]*kernel[7]+tmp[4055]*kernel[8];
				ans[3955]<=tmp[3854]*kernel[0]+tmp[3855]*kernel[1]+tmp[3856]*kernel[2]+tmp[3954]*kernel[3]+tmp[3955]*kernel[4]+tmp[3956]*kernel[5]+tmp[4054]*kernel[6]+tmp[4055]*kernel[7]+tmp[4056]*kernel[8];
				ans[3956]<=tmp[3855]*kernel[0]+tmp[3856]*kernel[1]+tmp[3857]*kernel[2]+tmp[3955]*kernel[3]+tmp[3956]*kernel[4]+tmp[3957]*kernel[5]+tmp[4055]*kernel[6]+tmp[4056]*kernel[7]+tmp[4057]*kernel[8];
				ans[3957]<=tmp[3856]*kernel[0]+tmp[3857]*kernel[1]+tmp[3858]*kernel[2]+tmp[3956]*kernel[3]+tmp[3957]*kernel[4]+tmp[3958]*kernel[5]+tmp[4056]*kernel[6]+tmp[4057]*kernel[7]+tmp[4058]*kernel[8];
				ans[3958]<=tmp[3857]*kernel[0]+tmp[3858]*kernel[1]+tmp[3859]*kernel[2]+tmp[3957]*kernel[3]+tmp[3958]*kernel[4]+tmp[3959]*kernel[5]+tmp[4057]*kernel[6]+tmp[4058]*kernel[7]+tmp[4059]*kernel[8];
				ans[3959]<=tmp[3858]*kernel[0]+tmp[3859]*kernel[1]+tmp[3860]*kernel[2]+tmp[3958]*kernel[3]+tmp[3959]*kernel[4]+tmp[3960]*kernel[5]+tmp[4058]*kernel[6]+tmp[4059]*kernel[7]+tmp[4060]*kernel[8];
				ans[3960]<=tmp[3859]*kernel[0]+tmp[3860]*kernel[1]+tmp[3861]*kernel[2]+tmp[3959]*kernel[3]+tmp[3960]*kernel[4]+tmp[3961]*kernel[5]+tmp[4059]*kernel[6]+tmp[4060]*kernel[7]+tmp[4061]*kernel[8];
				ans[3961]<=tmp[3860]*kernel[0]+tmp[3861]*kernel[1]+tmp[3862]*kernel[2]+tmp[3960]*kernel[3]+tmp[3961]*kernel[4]+tmp[3962]*kernel[5]+tmp[4060]*kernel[6]+tmp[4061]*kernel[7]+tmp[4062]*kernel[8];
				ans[3962]<=tmp[3861]*kernel[0]+tmp[3862]*kernel[1]+tmp[3863]*kernel[2]+tmp[3961]*kernel[3]+tmp[3962]*kernel[4]+tmp[3963]*kernel[5]+tmp[4061]*kernel[6]+tmp[4062]*kernel[7]+tmp[4063]*kernel[8];
				ans[3963]<=tmp[3862]*kernel[0]+tmp[3863]*kernel[1]+tmp[3864]*kernel[2]+tmp[3962]*kernel[3]+tmp[3963]*kernel[4]+tmp[3964]*kernel[5]+tmp[4062]*kernel[6]+tmp[4063]*kernel[7]+tmp[4064]*kernel[8];
				ans[3964]<=tmp[3863]*kernel[0]+tmp[3864]*kernel[1]+tmp[3865]*kernel[2]+tmp[3963]*kernel[3]+tmp[3964]*kernel[4]+tmp[3965]*kernel[5]+tmp[4063]*kernel[6]+tmp[4064]*kernel[7]+tmp[4065]*kernel[8];
				ans[3965]<=tmp[3864]*kernel[0]+tmp[3865]*kernel[1]+tmp[3866]*kernel[2]+tmp[3964]*kernel[3]+tmp[3965]*kernel[4]+tmp[3966]*kernel[5]+tmp[4064]*kernel[6]+tmp[4065]*kernel[7]+tmp[4066]*kernel[8];
				ans[3966]<=tmp[3865]*kernel[0]+tmp[3866]*kernel[1]+tmp[3867]*kernel[2]+tmp[3965]*kernel[3]+tmp[3966]*kernel[4]+tmp[3967]*kernel[5]+tmp[4065]*kernel[6]+tmp[4066]*kernel[7]+tmp[4067]*kernel[8];
				ans[3967]<=tmp[3866]*kernel[0]+tmp[3867]*kernel[1]+tmp[3868]*kernel[2]+tmp[3966]*kernel[3]+tmp[3967]*kernel[4]+tmp[3968]*kernel[5]+tmp[4066]*kernel[6]+tmp[4067]*kernel[7]+tmp[4068]*kernel[8];
				ans[3968]<=tmp[3867]*kernel[0]+tmp[3868]*kernel[1]+tmp[3869]*kernel[2]+tmp[3967]*kernel[3]+tmp[3968]*kernel[4]+tmp[3969]*kernel[5]+tmp[4067]*kernel[6]+tmp[4068]*kernel[7]+tmp[4069]*kernel[8];
				ans[3969]<=tmp[3868]*kernel[0]+tmp[3869]*kernel[1]+tmp[3870]*kernel[2]+tmp[3968]*kernel[3]+tmp[3969]*kernel[4]+tmp[3970]*kernel[5]+tmp[4068]*kernel[6]+tmp[4069]*kernel[7]+tmp[4070]*kernel[8];
				ans[3970]<=tmp[3869]*kernel[0]+tmp[3870]*kernel[1]+tmp[3871]*kernel[2]+tmp[3969]*kernel[3]+tmp[3970]*kernel[4]+tmp[3971]*kernel[5]+tmp[4069]*kernel[6]+tmp[4070]*kernel[7]+tmp[4071]*kernel[8];
				ans[3971]<=tmp[3870]*kernel[0]+tmp[3871]*kernel[1]+tmp[3872]*kernel[2]+tmp[3970]*kernel[3]+tmp[3971]*kernel[4]+tmp[3972]*kernel[5]+tmp[4070]*kernel[6]+tmp[4071]*kernel[7]+tmp[4072]*kernel[8];
				ans[3972]<=tmp[3871]*kernel[0]+tmp[3872]*kernel[1]+tmp[3873]*kernel[2]+tmp[3971]*kernel[3]+tmp[3972]*kernel[4]+tmp[3973]*kernel[5]+tmp[4071]*kernel[6]+tmp[4072]*kernel[7]+tmp[4073]*kernel[8];
				ans[3973]<=tmp[3872]*kernel[0]+tmp[3873]*kernel[1]+tmp[3874]*kernel[2]+tmp[3972]*kernel[3]+tmp[3973]*kernel[4]+tmp[3974]*kernel[5]+tmp[4072]*kernel[6]+tmp[4073]*kernel[7]+tmp[4074]*kernel[8];
				ans[3974]<=tmp[3873]*kernel[0]+tmp[3874]*kernel[1]+tmp[3875]*kernel[2]+tmp[3973]*kernel[3]+tmp[3974]*kernel[4]+tmp[3975]*kernel[5]+tmp[4073]*kernel[6]+tmp[4074]*kernel[7]+tmp[4075]*kernel[8];
				ans[3975]<=tmp[3874]*kernel[0]+tmp[3875]*kernel[1]+tmp[3876]*kernel[2]+tmp[3974]*kernel[3]+tmp[3975]*kernel[4]+tmp[3976]*kernel[5]+tmp[4074]*kernel[6]+tmp[4075]*kernel[7]+tmp[4076]*kernel[8];
				ans[3976]<=tmp[3875]*kernel[0]+tmp[3876]*kernel[1]+tmp[3877]*kernel[2]+tmp[3975]*kernel[3]+tmp[3976]*kernel[4]+tmp[3977]*kernel[5]+tmp[4075]*kernel[6]+tmp[4076]*kernel[7]+tmp[4077]*kernel[8];
				ans[3977]<=tmp[3876]*kernel[0]+tmp[3877]*kernel[1]+tmp[3878]*kernel[2]+tmp[3976]*kernel[3]+tmp[3977]*kernel[4]+tmp[3978]*kernel[5]+tmp[4076]*kernel[6]+tmp[4077]*kernel[7]+tmp[4078]*kernel[8];
				ans[3978]<=tmp[3877]*kernel[0]+tmp[3878]*kernel[1]+tmp[3879]*kernel[2]+tmp[3977]*kernel[3]+tmp[3978]*kernel[4]+tmp[3979]*kernel[5]+tmp[4077]*kernel[6]+tmp[4078]*kernel[7]+tmp[4079]*kernel[8];
				ans[3979]<=tmp[3878]*kernel[0]+tmp[3879]*kernel[1]+tmp[3880]*kernel[2]+tmp[3978]*kernel[3]+tmp[3979]*kernel[4]+tmp[3980]*kernel[5]+tmp[4078]*kernel[6]+tmp[4079]*kernel[7]+tmp[4080]*kernel[8];
				ans[3980]<=tmp[3879]*kernel[0]+tmp[3880]*kernel[1]+tmp[3881]*kernel[2]+tmp[3979]*kernel[3]+tmp[3980]*kernel[4]+tmp[3981]*kernel[5]+tmp[4079]*kernel[6]+tmp[4080]*kernel[7]+tmp[4081]*kernel[8];
				ans[3981]<=tmp[3880]*kernel[0]+tmp[3881]*kernel[1]+tmp[3882]*kernel[2]+tmp[3980]*kernel[3]+tmp[3981]*kernel[4]+tmp[3982]*kernel[5]+tmp[4080]*kernel[6]+tmp[4081]*kernel[7]+tmp[4082]*kernel[8];
				ans[3982]<=tmp[3881]*kernel[0]+tmp[3882]*kernel[1]+tmp[3883]*kernel[2]+tmp[3981]*kernel[3]+tmp[3982]*kernel[4]+tmp[3983]*kernel[5]+tmp[4081]*kernel[6]+tmp[4082]*kernel[7]+tmp[4083]*kernel[8];
				ans[3983]<=tmp[3882]*kernel[0]+tmp[3883]*kernel[1]+tmp[3884]*kernel[2]+tmp[3982]*kernel[3]+tmp[3983]*kernel[4]+tmp[3984]*kernel[5]+tmp[4082]*kernel[6]+tmp[4083]*kernel[7]+tmp[4084]*kernel[8];
				ans[3984]<=tmp[3883]*kernel[0]+tmp[3884]*kernel[1]+tmp[3885]*kernel[2]+tmp[3983]*kernel[3]+tmp[3984]*kernel[4]+tmp[3985]*kernel[5]+tmp[4083]*kernel[6]+tmp[4084]*kernel[7]+tmp[4085]*kernel[8];
				ans[3985]<=tmp[3884]*kernel[0]+tmp[3885]*kernel[1]+tmp[3886]*kernel[2]+tmp[3984]*kernel[3]+tmp[3985]*kernel[4]+tmp[3986]*kernel[5]+tmp[4084]*kernel[6]+tmp[4085]*kernel[7]+tmp[4086]*kernel[8];
				ans[3986]<=tmp[3885]*kernel[0]+tmp[3886]*kernel[1]+tmp[3887]*kernel[2]+tmp[3985]*kernel[3]+tmp[3986]*kernel[4]+tmp[3987]*kernel[5]+tmp[4085]*kernel[6]+tmp[4086]*kernel[7]+tmp[4087]*kernel[8];
				ans[3987]<=tmp[3886]*kernel[0]+tmp[3887]*kernel[1]+tmp[3888]*kernel[2]+tmp[3986]*kernel[3]+tmp[3987]*kernel[4]+tmp[3988]*kernel[5]+tmp[4086]*kernel[6]+tmp[4087]*kernel[7]+tmp[4088]*kernel[8];
				ans[3988]<=tmp[3887]*kernel[0]+tmp[3888]*kernel[1]+tmp[3889]*kernel[2]+tmp[3987]*kernel[3]+tmp[3988]*kernel[4]+tmp[3989]*kernel[5]+tmp[4087]*kernel[6]+tmp[4088]*kernel[7]+tmp[4089]*kernel[8];
				ans[3989]<=tmp[3888]*kernel[0]+tmp[3889]*kernel[1]+tmp[3890]*kernel[2]+tmp[3988]*kernel[3]+tmp[3989]*kernel[4]+tmp[3990]*kernel[5]+tmp[4088]*kernel[6]+tmp[4089]*kernel[7]+tmp[4090]*kernel[8];
				ans[3990]<=tmp[3889]*kernel[0]+tmp[3890]*kernel[1]+tmp[3891]*kernel[2]+tmp[3989]*kernel[3]+tmp[3990]*kernel[4]+tmp[3991]*kernel[5]+tmp[4089]*kernel[6]+tmp[4090]*kernel[7]+tmp[4091]*kernel[8];
				ans[3991]<=tmp[3890]*kernel[0]+tmp[3891]*kernel[1]+tmp[3892]*kernel[2]+tmp[3990]*kernel[3]+tmp[3991]*kernel[4]+tmp[3992]*kernel[5]+tmp[4090]*kernel[6]+tmp[4091]*kernel[7]+tmp[4092]*kernel[8];
				ans[3992]<=tmp[3891]*kernel[0]+tmp[3892]*kernel[1]+tmp[3893]*kernel[2]+tmp[3991]*kernel[3]+tmp[3992]*kernel[4]+tmp[3993]*kernel[5]+tmp[4091]*kernel[6]+tmp[4092]*kernel[7]+tmp[4093]*kernel[8];
				ans[3993]<=tmp[3892]*kernel[0]+tmp[3893]*kernel[1]+tmp[3894]*kernel[2]+tmp[3992]*kernel[3]+tmp[3993]*kernel[4]+tmp[3994]*kernel[5]+tmp[4092]*kernel[6]+tmp[4093]*kernel[7]+tmp[4094]*kernel[8];
				ans[3994]<=tmp[3893]*kernel[0]+tmp[3894]*kernel[1]+tmp[3895]*kernel[2]+tmp[3993]*kernel[3]+tmp[3994]*kernel[4]+tmp[3995]*kernel[5]+tmp[4093]*kernel[6]+tmp[4094]*kernel[7]+tmp[4095]*kernel[8];
				ans[3995]<=tmp[3894]*kernel[0]+tmp[3895]*kernel[1]+tmp[3896]*kernel[2]+tmp[3994]*kernel[3]+tmp[3995]*kernel[4]+tmp[3996]*kernel[5]+tmp[4094]*kernel[6]+tmp[4095]*kernel[7]+tmp[4096]*kernel[8];
				ans[3996]<=tmp[3895]*kernel[0]+tmp[3896]*kernel[1]+tmp[3897]*kernel[2]+tmp[3995]*kernel[3]+tmp[3996]*kernel[4]+tmp[3997]*kernel[5]+tmp[4095]*kernel[6]+tmp[4096]*kernel[7]+tmp[4097]*kernel[8];
				ans[3997]<=tmp[3896]*kernel[0]+tmp[3897]*kernel[1]+tmp[3898]*kernel[2]+tmp[3996]*kernel[3]+tmp[3997]*kernel[4]+tmp[3998]*kernel[5]+tmp[4096]*kernel[6]+tmp[4097]*kernel[7]+tmp[4098]*kernel[8];
				ans[3998]<=tmp[3897]*kernel[0]+tmp[3898]*kernel[1]+tmp[3899]*kernel[2]+tmp[3997]*kernel[3]+tmp[3998]*kernel[4]+tmp[3999]*kernel[5]+tmp[4097]*kernel[6]+tmp[4098]*kernel[7]+tmp[4099]*kernel[8];
				ans[3999]<=tmp[3898]*kernel[0]+tmp[3899]*kernel[1]+tmp[3998]*kernel[3]+tmp[3999]*kernel[4]+tmp[4098]*kernel[6]+tmp[4099]*kernel[7];
				ans[4000]<=tmp[3900]*kernel[1]+tmp[3901]*kernel[2]+tmp[4000]*kernel[4]+tmp[4001]*kernel[5]+tmp[4100]*kernel[7]+tmp[4101]*kernel[8];
				ans[4001]<=tmp[3900]*kernel[0]+tmp[3901]*kernel[1]+tmp[3902]*kernel[2]+tmp[4000]*kernel[3]+tmp[4001]*kernel[4]+tmp[4002]*kernel[5]+tmp[4100]*kernel[6]+tmp[4101]*kernel[7]+tmp[4102]*kernel[8];
				ans[4002]<=tmp[3901]*kernel[0]+tmp[3902]*kernel[1]+tmp[3903]*kernel[2]+tmp[4001]*kernel[3]+tmp[4002]*kernel[4]+tmp[4003]*kernel[5]+tmp[4101]*kernel[6]+tmp[4102]*kernel[7]+tmp[4103]*kernel[8];
				ans[4003]<=tmp[3902]*kernel[0]+tmp[3903]*kernel[1]+tmp[3904]*kernel[2]+tmp[4002]*kernel[3]+tmp[4003]*kernel[4]+tmp[4004]*kernel[5]+tmp[4102]*kernel[6]+tmp[4103]*kernel[7]+tmp[4104]*kernel[8];
				ans[4004]<=tmp[3903]*kernel[0]+tmp[3904]*kernel[1]+tmp[3905]*kernel[2]+tmp[4003]*kernel[3]+tmp[4004]*kernel[4]+tmp[4005]*kernel[5]+tmp[4103]*kernel[6]+tmp[4104]*kernel[7]+tmp[4105]*kernel[8];
				ans[4005]<=tmp[3904]*kernel[0]+tmp[3905]*kernel[1]+tmp[3906]*kernel[2]+tmp[4004]*kernel[3]+tmp[4005]*kernel[4]+tmp[4006]*kernel[5]+tmp[4104]*kernel[6]+tmp[4105]*kernel[7]+tmp[4106]*kernel[8];
				ans[4006]<=tmp[3905]*kernel[0]+tmp[3906]*kernel[1]+tmp[3907]*kernel[2]+tmp[4005]*kernel[3]+tmp[4006]*kernel[4]+tmp[4007]*kernel[5]+tmp[4105]*kernel[6]+tmp[4106]*kernel[7]+tmp[4107]*kernel[8];
				ans[4007]<=tmp[3906]*kernel[0]+tmp[3907]*kernel[1]+tmp[3908]*kernel[2]+tmp[4006]*kernel[3]+tmp[4007]*kernel[4]+tmp[4008]*kernel[5]+tmp[4106]*kernel[6]+tmp[4107]*kernel[7]+tmp[4108]*kernel[8];
				ans[4008]<=tmp[3907]*kernel[0]+tmp[3908]*kernel[1]+tmp[3909]*kernel[2]+tmp[4007]*kernel[3]+tmp[4008]*kernel[4]+tmp[4009]*kernel[5]+tmp[4107]*kernel[6]+tmp[4108]*kernel[7]+tmp[4109]*kernel[8];
				ans[4009]<=tmp[3908]*kernel[0]+tmp[3909]*kernel[1]+tmp[3910]*kernel[2]+tmp[4008]*kernel[3]+tmp[4009]*kernel[4]+tmp[4010]*kernel[5]+tmp[4108]*kernel[6]+tmp[4109]*kernel[7]+tmp[4110]*kernel[8];
				ans[4010]<=tmp[3909]*kernel[0]+tmp[3910]*kernel[1]+tmp[3911]*kernel[2]+tmp[4009]*kernel[3]+tmp[4010]*kernel[4]+tmp[4011]*kernel[5]+tmp[4109]*kernel[6]+tmp[4110]*kernel[7]+tmp[4111]*kernel[8];
				ans[4011]<=tmp[3910]*kernel[0]+tmp[3911]*kernel[1]+tmp[3912]*kernel[2]+tmp[4010]*kernel[3]+tmp[4011]*kernel[4]+tmp[4012]*kernel[5]+tmp[4110]*kernel[6]+tmp[4111]*kernel[7]+tmp[4112]*kernel[8];
				ans[4012]<=tmp[3911]*kernel[0]+tmp[3912]*kernel[1]+tmp[3913]*kernel[2]+tmp[4011]*kernel[3]+tmp[4012]*kernel[4]+tmp[4013]*kernel[5]+tmp[4111]*kernel[6]+tmp[4112]*kernel[7]+tmp[4113]*kernel[8];
				ans[4013]<=tmp[3912]*kernel[0]+tmp[3913]*kernel[1]+tmp[3914]*kernel[2]+tmp[4012]*kernel[3]+tmp[4013]*kernel[4]+tmp[4014]*kernel[5]+tmp[4112]*kernel[6]+tmp[4113]*kernel[7]+tmp[4114]*kernel[8];
				ans[4014]<=tmp[3913]*kernel[0]+tmp[3914]*kernel[1]+tmp[3915]*kernel[2]+tmp[4013]*kernel[3]+tmp[4014]*kernel[4]+tmp[4015]*kernel[5]+tmp[4113]*kernel[6]+tmp[4114]*kernel[7]+tmp[4115]*kernel[8];
				ans[4015]<=tmp[3914]*kernel[0]+tmp[3915]*kernel[1]+tmp[3916]*kernel[2]+tmp[4014]*kernel[3]+tmp[4015]*kernel[4]+tmp[4016]*kernel[5]+tmp[4114]*kernel[6]+tmp[4115]*kernel[7]+tmp[4116]*kernel[8];
				ans[4016]<=tmp[3915]*kernel[0]+tmp[3916]*kernel[1]+tmp[3917]*kernel[2]+tmp[4015]*kernel[3]+tmp[4016]*kernel[4]+tmp[4017]*kernel[5]+tmp[4115]*kernel[6]+tmp[4116]*kernel[7]+tmp[4117]*kernel[8];
				ans[4017]<=tmp[3916]*kernel[0]+tmp[3917]*kernel[1]+tmp[3918]*kernel[2]+tmp[4016]*kernel[3]+tmp[4017]*kernel[4]+tmp[4018]*kernel[5]+tmp[4116]*kernel[6]+tmp[4117]*kernel[7]+tmp[4118]*kernel[8];
				ans[4018]<=tmp[3917]*kernel[0]+tmp[3918]*kernel[1]+tmp[3919]*kernel[2]+tmp[4017]*kernel[3]+tmp[4018]*kernel[4]+tmp[4019]*kernel[5]+tmp[4117]*kernel[6]+tmp[4118]*kernel[7]+tmp[4119]*kernel[8];
				ans[4019]<=tmp[3918]*kernel[0]+tmp[3919]*kernel[1]+tmp[3920]*kernel[2]+tmp[4018]*kernel[3]+tmp[4019]*kernel[4]+tmp[4020]*kernel[5]+tmp[4118]*kernel[6]+tmp[4119]*kernel[7]+tmp[4120]*kernel[8];
				ans[4020]<=tmp[3919]*kernel[0]+tmp[3920]*kernel[1]+tmp[3921]*kernel[2]+tmp[4019]*kernel[3]+tmp[4020]*kernel[4]+tmp[4021]*kernel[5]+tmp[4119]*kernel[6]+tmp[4120]*kernel[7]+tmp[4121]*kernel[8];
				ans[4021]<=tmp[3920]*kernel[0]+tmp[3921]*kernel[1]+tmp[3922]*kernel[2]+tmp[4020]*kernel[3]+tmp[4021]*kernel[4]+tmp[4022]*kernel[5]+tmp[4120]*kernel[6]+tmp[4121]*kernel[7]+tmp[4122]*kernel[8];
				ans[4022]<=tmp[3921]*kernel[0]+tmp[3922]*kernel[1]+tmp[3923]*kernel[2]+tmp[4021]*kernel[3]+tmp[4022]*kernel[4]+tmp[4023]*kernel[5]+tmp[4121]*kernel[6]+tmp[4122]*kernel[7]+tmp[4123]*kernel[8];
				ans[4023]<=tmp[3922]*kernel[0]+tmp[3923]*kernel[1]+tmp[3924]*kernel[2]+tmp[4022]*kernel[3]+tmp[4023]*kernel[4]+tmp[4024]*kernel[5]+tmp[4122]*kernel[6]+tmp[4123]*kernel[7]+tmp[4124]*kernel[8];
				ans[4024]<=tmp[3923]*kernel[0]+tmp[3924]*kernel[1]+tmp[3925]*kernel[2]+tmp[4023]*kernel[3]+tmp[4024]*kernel[4]+tmp[4025]*kernel[5]+tmp[4123]*kernel[6]+tmp[4124]*kernel[7]+tmp[4125]*kernel[8];
				ans[4025]<=tmp[3924]*kernel[0]+tmp[3925]*kernel[1]+tmp[3926]*kernel[2]+tmp[4024]*kernel[3]+tmp[4025]*kernel[4]+tmp[4026]*kernel[5]+tmp[4124]*kernel[6]+tmp[4125]*kernel[7]+tmp[4126]*kernel[8];
				ans[4026]<=tmp[3925]*kernel[0]+tmp[3926]*kernel[1]+tmp[3927]*kernel[2]+tmp[4025]*kernel[3]+tmp[4026]*kernel[4]+tmp[4027]*kernel[5]+tmp[4125]*kernel[6]+tmp[4126]*kernel[7]+tmp[4127]*kernel[8];
				ans[4027]<=tmp[3926]*kernel[0]+tmp[3927]*kernel[1]+tmp[3928]*kernel[2]+tmp[4026]*kernel[3]+tmp[4027]*kernel[4]+tmp[4028]*kernel[5]+tmp[4126]*kernel[6]+tmp[4127]*kernel[7]+tmp[4128]*kernel[8];
				ans[4028]<=tmp[3927]*kernel[0]+tmp[3928]*kernel[1]+tmp[3929]*kernel[2]+tmp[4027]*kernel[3]+tmp[4028]*kernel[4]+tmp[4029]*kernel[5]+tmp[4127]*kernel[6]+tmp[4128]*kernel[7]+tmp[4129]*kernel[8];
				ans[4029]<=tmp[3928]*kernel[0]+tmp[3929]*kernel[1]+tmp[3930]*kernel[2]+tmp[4028]*kernel[3]+tmp[4029]*kernel[4]+tmp[4030]*kernel[5]+tmp[4128]*kernel[6]+tmp[4129]*kernel[7]+tmp[4130]*kernel[8];
				ans[4030]<=tmp[3929]*kernel[0]+tmp[3930]*kernel[1]+tmp[3931]*kernel[2]+tmp[4029]*kernel[3]+tmp[4030]*kernel[4]+tmp[4031]*kernel[5]+tmp[4129]*kernel[6]+tmp[4130]*kernel[7]+tmp[4131]*kernel[8];
				ans[4031]<=tmp[3930]*kernel[0]+tmp[3931]*kernel[1]+tmp[3932]*kernel[2]+tmp[4030]*kernel[3]+tmp[4031]*kernel[4]+tmp[4032]*kernel[5]+tmp[4130]*kernel[6]+tmp[4131]*kernel[7]+tmp[4132]*kernel[8];
				ans[4032]<=tmp[3931]*kernel[0]+tmp[3932]*kernel[1]+tmp[3933]*kernel[2]+tmp[4031]*kernel[3]+tmp[4032]*kernel[4]+tmp[4033]*kernel[5]+tmp[4131]*kernel[6]+tmp[4132]*kernel[7]+tmp[4133]*kernel[8];
				ans[4033]<=tmp[3932]*kernel[0]+tmp[3933]*kernel[1]+tmp[3934]*kernel[2]+tmp[4032]*kernel[3]+tmp[4033]*kernel[4]+tmp[4034]*kernel[5]+tmp[4132]*kernel[6]+tmp[4133]*kernel[7]+tmp[4134]*kernel[8];
				ans[4034]<=tmp[3933]*kernel[0]+tmp[3934]*kernel[1]+tmp[3935]*kernel[2]+tmp[4033]*kernel[3]+tmp[4034]*kernel[4]+tmp[4035]*kernel[5]+tmp[4133]*kernel[6]+tmp[4134]*kernel[7]+tmp[4135]*kernel[8];
				ans[4035]<=tmp[3934]*kernel[0]+tmp[3935]*kernel[1]+tmp[3936]*kernel[2]+tmp[4034]*kernel[3]+tmp[4035]*kernel[4]+tmp[4036]*kernel[5]+tmp[4134]*kernel[6]+tmp[4135]*kernel[7]+tmp[4136]*kernel[8];
				ans[4036]<=tmp[3935]*kernel[0]+tmp[3936]*kernel[1]+tmp[3937]*kernel[2]+tmp[4035]*kernel[3]+tmp[4036]*kernel[4]+tmp[4037]*kernel[5]+tmp[4135]*kernel[6]+tmp[4136]*kernel[7]+tmp[4137]*kernel[8];
				ans[4037]<=tmp[3936]*kernel[0]+tmp[3937]*kernel[1]+tmp[3938]*kernel[2]+tmp[4036]*kernel[3]+tmp[4037]*kernel[4]+tmp[4038]*kernel[5]+tmp[4136]*kernel[6]+tmp[4137]*kernel[7]+tmp[4138]*kernel[8];
				ans[4038]<=tmp[3937]*kernel[0]+tmp[3938]*kernel[1]+tmp[3939]*kernel[2]+tmp[4037]*kernel[3]+tmp[4038]*kernel[4]+tmp[4039]*kernel[5]+tmp[4137]*kernel[6]+tmp[4138]*kernel[7]+tmp[4139]*kernel[8];
				ans[4039]<=tmp[3938]*kernel[0]+tmp[3939]*kernel[1]+tmp[3940]*kernel[2]+tmp[4038]*kernel[3]+tmp[4039]*kernel[4]+tmp[4040]*kernel[5]+tmp[4138]*kernel[6]+tmp[4139]*kernel[7]+tmp[4140]*kernel[8];
				ans[4040]<=tmp[3939]*kernel[0]+tmp[3940]*kernel[1]+tmp[3941]*kernel[2]+tmp[4039]*kernel[3]+tmp[4040]*kernel[4]+tmp[4041]*kernel[5]+tmp[4139]*kernel[6]+tmp[4140]*kernel[7]+tmp[4141]*kernel[8];
				ans[4041]<=tmp[3940]*kernel[0]+tmp[3941]*kernel[1]+tmp[3942]*kernel[2]+tmp[4040]*kernel[3]+tmp[4041]*kernel[4]+tmp[4042]*kernel[5]+tmp[4140]*kernel[6]+tmp[4141]*kernel[7]+tmp[4142]*kernel[8];
				ans[4042]<=tmp[3941]*kernel[0]+tmp[3942]*kernel[1]+tmp[3943]*kernel[2]+tmp[4041]*kernel[3]+tmp[4042]*kernel[4]+tmp[4043]*kernel[5]+tmp[4141]*kernel[6]+tmp[4142]*kernel[7]+tmp[4143]*kernel[8];
				ans[4043]<=tmp[3942]*kernel[0]+tmp[3943]*kernel[1]+tmp[3944]*kernel[2]+tmp[4042]*kernel[3]+tmp[4043]*kernel[4]+tmp[4044]*kernel[5]+tmp[4142]*kernel[6]+tmp[4143]*kernel[7]+tmp[4144]*kernel[8];
				ans[4044]<=tmp[3943]*kernel[0]+tmp[3944]*kernel[1]+tmp[3945]*kernel[2]+tmp[4043]*kernel[3]+tmp[4044]*kernel[4]+tmp[4045]*kernel[5]+tmp[4143]*kernel[6]+tmp[4144]*kernel[7]+tmp[4145]*kernel[8];
				ans[4045]<=tmp[3944]*kernel[0]+tmp[3945]*kernel[1]+tmp[3946]*kernel[2]+tmp[4044]*kernel[3]+tmp[4045]*kernel[4]+tmp[4046]*kernel[5]+tmp[4144]*kernel[6]+tmp[4145]*kernel[7]+tmp[4146]*kernel[8];
				ans[4046]<=tmp[3945]*kernel[0]+tmp[3946]*kernel[1]+tmp[3947]*kernel[2]+tmp[4045]*kernel[3]+tmp[4046]*kernel[4]+tmp[4047]*kernel[5]+tmp[4145]*kernel[6]+tmp[4146]*kernel[7]+tmp[4147]*kernel[8];
				ans[4047]<=tmp[3946]*kernel[0]+tmp[3947]*kernel[1]+tmp[3948]*kernel[2]+tmp[4046]*kernel[3]+tmp[4047]*kernel[4]+tmp[4048]*kernel[5]+tmp[4146]*kernel[6]+tmp[4147]*kernel[7]+tmp[4148]*kernel[8];
				ans[4048]<=tmp[3947]*kernel[0]+tmp[3948]*kernel[1]+tmp[3949]*kernel[2]+tmp[4047]*kernel[3]+tmp[4048]*kernel[4]+tmp[4049]*kernel[5]+tmp[4147]*kernel[6]+tmp[4148]*kernel[7]+tmp[4149]*kernel[8];
				ans[4049]<=tmp[3948]*kernel[0]+tmp[3949]*kernel[1]+tmp[3950]*kernel[2]+tmp[4048]*kernel[3]+tmp[4049]*kernel[4]+tmp[4050]*kernel[5]+tmp[4148]*kernel[6]+tmp[4149]*kernel[7]+tmp[4150]*kernel[8];
				ans[4050]<=tmp[3949]*kernel[0]+tmp[3950]*kernel[1]+tmp[3951]*kernel[2]+tmp[4049]*kernel[3]+tmp[4050]*kernel[4]+tmp[4051]*kernel[5]+tmp[4149]*kernel[6]+tmp[4150]*kernel[7]+tmp[4151]*kernel[8];
				ans[4051]<=tmp[3950]*kernel[0]+tmp[3951]*kernel[1]+tmp[3952]*kernel[2]+tmp[4050]*kernel[3]+tmp[4051]*kernel[4]+tmp[4052]*kernel[5]+tmp[4150]*kernel[6]+tmp[4151]*kernel[7]+tmp[4152]*kernel[8];
				ans[4052]<=tmp[3951]*kernel[0]+tmp[3952]*kernel[1]+tmp[3953]*kernel[2]+tmp[4051]*kernel[3]+tmp[4052]*kernel[4]+tmp[4053]*kernel[5]+tmp[4151]*kernel[6]+tmp[4152]*kernel[7]+tmp[4153]*kernel[8];
				ans[4053]<=tmp[3952]*kernel[0]+tmp[3953]*kernel[1]+tmp[3954]*kernel[2]+tmp[4052]*kernel[3]+tmp[4053]*kernel[4]+tmp[4054]*kernel[5]+tmp[4152]*kernel[6]+tmp[4153]*kernel[7]+tmp[4154]*kernel[8];
				ans[4054]<=tmp[3953]*kernel[0]+tmp[3954]*kernel[1]+tmp[3955]*kernel[2]+tmp[4053]*kernel[3]+tmp[4054]*kernel[4]+tmp[4055]*kernel[5]+tmp[4153]*kernel[6]+tmp[4154]*kernel[7]+tmp[4155]*kernel[8];
				ans[4055]<=tmp[3954]*kernel[0]+tmp[3955]*kernel[1]+tmp[3956]*kernel[2]+tmp[4054]*kernel[3]+tmp[4055]*kernel[4]+tmp[4056]*kernel[5]+tmp[4154]*kernel[6]+tmp[4155]*kernel[7]+tmp[4156]*kernel[8];
				ans[4056]<=tmp[3955]*kernel[0]+tmp[3956]*kernel[1]+tmp[3957]*kernel[2]+tmp[4055]*kernel[3]+tmp[4056]*kernel[4]+tmp[4057]*kernel[5]+tmp[4155]*kernel[6]+tmp[4156]*kernel[7]+tmp[4157]*kernel[8];
				ans[4057]<=tmp[3956]*kernel[0]+tmp[3957]*kernel[1]+tmp[3958]*kernel[2]+tmp[4056]*kernel[3]+tmp[4057]*kernel[4]+tmp[4058]*kernel[5]+tmp[4156]*kernel[6]+tmp[4157]*kernel[7]+tmp[4158]*kernel[8];
				ans[4058]<=tmp[3957]*kernel[0]+tmp[3958]*kernel[1]+tmp[3959]*kernel[2]+tmp[4057]*kernel[3]+tmp[4058]*kernel[4]+tmp[4059]*kernel[5]+tmp[4157]*kernel[6]+tmp[4158]*kernel[7]+tmp[4159]*kernel[8];
				ans[4059]<=tmp[3958]*kernel[0]+tmp[3959]*kernel[1]+tmp[3960]*kernel[2]+tmp[4058]*kernel[3]+tmp[4059]*kernel[4]+tmp[4060]*kernel[5]+tmp[4158]*kernel[6]+tmp[4159]*kernel[7]+tmp[4160]*kernel[8];
				ans[4060]<=tmp[3959]*kernel[0]+tmp[3960]*kernel[1]+tmp[3961]*kernel[2]+tmp[4059]*kernel[3]+tmp[4060]*kernel[4]+tmp[4061]*kernel[5]+tmp[4159]*kernel[6]+tmp[4160]*kernel[7]+tmp[4161]*kernel[8];
				ans[4061]<=tmp[3960]*kernel[0]+tmp[3961]*kernel[1]+tmp[3962]*kernel[2]+tmp[4060]*kernel[3]+tmp[4061]*kernel[4]+tmp[4062]*kernel[5]+tmp[4160]*kernel[6]+tmp[4161]*kernel[7]+tmp[4162]*kernel[8];
				ans[4062]<=tmp[3961]*kernel[0]+tmp[3962]*kernel[1]+tmp[3963]*kernel[2]+tmp[4061]*kernel[3]+tmp[4062]*kernel[4]+tmp[4063]*kernel[5]+tmp[4161]*kernel[6]+tmp[4162]*kernel[7]+tmp[4163]*kernel[8];
				ans[4063]<=tmp[3962]*kernel[0]+tmp[3963]*kernel[1]+tmp[3964]*kernel[2]+tmp[4062]*kernel[3]+tmp[4063]*kernel[4]+tmp[4064]*kernel[5]+tmp[4162]*kernel[6]+tmp[4163]*kernel[7]+tmp[4164]*kernel[8];
				ans[4064]<=tmp[3963]*kernel[0]+tmp[3964]*kernel[1]+tmp[3965]*kernel[2]+tmp[4063]*kernel[3]+tmp[4064]*kernel[4]+tmp[4065]*kernel[5]+tmp[4163]*kernel[6]+tmp[4164]*kernel[7]+tmp[4165]*kernel[8];
				ans[4065]<=tmp[3964]*kernel[0]+tmp[3965]*kernel[1]+tmp[3966]*kernel[2]+tmp[4064]*kernel[3]+tmp[4065]*kernel[4]+tmp[4066]*kernel[5]+tmp[4164]*kernel[6]+tmp[4165]*kernel[7]+tmp[4166]*kernel[8];
				ans[4066]<=tmp[3965]*kernel[0]+tmp[3966]*kernel[1]+tmp[3967]*kernel[2]+tmp[4065]*kernel[3]+tmp[4066]*kernel[4]+tmp[4067]*kernel[5]+tmp[4165]*kernel[6]+tmp[4166]*kernel[7]+tmp[4167]*kernel[8];
				ans[4067]<=tmp[3966]*kernel[0]+tmp[3967]*kernel[1]+tmp[3968]*kernel[2]+tmp[4066]*kernel[3]+tmp[4067]*kernel[4]+tmp[4068]*kernel[5]+tmp[4166]*kernel[6]+tmp[4167]*kernel[7]+tmp[4168]*kernel[8];
				ans[4068]<=tmp[3967]*kernel[0]+tmp[3968]*kernel[1]+tmp[3969]*kernel[2]+tmp[4067]*kernel[3]+tmp[4068]*kernel[4]+tmp[4069]*kernel[5]+tmp[4167]*kernel[6]+tmp[4168]*kernel[7]+tmp[4169]*kernel[8];
				ans[4069]<=tmp[3968]*kernel[0]+tmp[3969]*kernel[1]+tmp[3970]*kernel[2]+tmp[4068]*kernel[3]+tmp[4069]*kernel[4]+tmp[4070]*kernel[5]+tmp[4168]*kernel[6]+tmp[4169]*kernel[7]+tmp[4170]*kernel[8];
				ans[4070]<=tmp[3969]*kernel[0]+tmp[3970]*kernel[1]+tmp[3971]*kernel[2]+tmp[4069]*kernel[3]+tmp[4070]*kernel[4]+tmp[4071]*kernel[5]+tmp[4169]*kernel[6]+tmp[4170]*kernel[7]+tmp[4171]*kernel[8];
				ans[4071]<=tmp[3970]*kernel[0]+tmp[3971]*kernel[1]+tmp[3972]*kernel[2]+tmp[4070]*kernel[3]+tmp[4071]*kernel[4]+tmp[4072]*kernel[5]+tmp[4170]*kernel[6]+tmp[4171]*kernel[7]+tmp[4172]*kernel[8];
				ans[4072]<=tmp[3971]*kernel[0]+tmp[3972]*kernel[1]+tmp[3973]*kernel[2]+tmp[4071]*kernel[3]+tmp[4072]*kernel[4]+tmp[4073]*kernel[5]+tmp[4171]*kernel[6]+tmp[4172]*kernel[7]+tmp[4173]*kernel[8];
				ans[4073]<=tmp[3972]*kernel[0]+tmp[3973]*kernel[1]+tmp[3974]*kernel[2]+tmp[4072]*kernel[3]+tmp[4073]*kernel[4]+tmp[4074]*kernel[5]+tmp[4172]*kernel[6]+tmp[4173]*kernel[7]+tmp[4174]*kernel[8];
				ans[4074]<=tmp[3973]*kernel[0]+tmp[3974]*kernel[1]+tmp[3975]*kernel[2]+tmp[4073]*kernel[3]+tmp[4074]*kernel[4]+tmp[4075]*kernel[5]+tmp[4173]*kernel[6]+tmp[4174]*kernel[7]+tmp[4175]*kernel[8];
				ans[4075]<=tmp[3974]*kernel[0]+tmp[3975]*kernel[1]+tmp[3976]*kernel[2]+tmp[4074]*kernel[3]+tmp[4075]*kernel[4]+tmp[4076]*kernel[5]+tmp[4174]*kernel[6]+tmp[4175]*kernel[7]+tmp[4176]*kernel[8];
				ans[4076]<=tmp[3975]*kernel[0]+tmp[3976]*kernel[1]+tmp[3977]*kernel[2]+tmp[4075]*kernel[3]+tmp[4076]*kernel[4]+tmp[4077]*kernel[5]+tmp[4175]*kernel[6]+tmp[4176]*kernel[7]+tmp[4177]*kernel[8];
				ans[4077]<=tmp[3976]*kernel[0]+tmp[3977]*kernel[1]+tmp[3978]*kernel[2]+tmp[4076]*kernel[3]+tmp[4077]*kernel[4]+tmp[4078]*kernel[5]+tmp[4176]*kernel[6]+tmp[4177]*kernel[7]+tmp[4178]*kernel[8];
				ans[4078]<=tmp[3977]*kernel[0]+tmp[3978]*kernel[1]+tmp[3979]*kernel[2]+tmp[4077]*kernel[3]+tmp[4078]*kernel[4]+tmp[4079]*kernel[5]+tmp[4177]*kernel[6]+tmp[4178]*kernel[7]+tmp[4179]*kernel[8];
				ans[4079]<=tmp[3978]*kernel[0]+tmp[3979]*kernel[1]+tmp[3980]*kernel[2]+tmp[4078]*kernel[3]+tmp[4079]*kernel[4]+tmp[4080]*kernel[5]+tmp[4178]*kernel[6]+tmp[4179]*kernel[7]+tmp[4180]*kernel[8];
				ans[4080]<=tmp[3979]*kernel[0]+tmp[3980]*kernel[1]+tmp[3981]*kernel[2]+tmp[4079]*kernel[3]+tmp[4080]*kernel[4]+tmp[4081]*kernel[5]+tmp[4179]*kernel[6]+tmp[4180]*kernel[7]+tmp[4181]*kernel[8];
				ans[4081]<=tmp[3980]*kernel[0]+tmp[3981]*kernel[1]+tmp[3982]*kernel[2]+tmp[4080]*kernel[3]+tmp[4081]*kernel[4]+tmp[4082]*kernel[5]+tmp[4180]*kernel[6]+tmp[4181]*kernel[7]+tmp[4182]*kernel[8];
				ans[4082]<=tmp[3981]*kernel[0]+tmp[3982]*kernel[1]+tmp[3983]*kernel[2]+tmp[4081]*kernel[3]+tmp[4082]*kernel[4]+tmp[4083]*kernel[5]+tmp[4181]*kernel[6]+tmp[4182]*kernel[7]+tmp[4183]*kernel[8];
				ans[4083]<=tmp[3982]*kernel[0]+tmp[3983]*kernel[1]+tmp[3984]*kernel[2]+tmp[4082]*kernel[3]+tmp[4083]*kernel[4]+tmp[4084]*kernel[5]+tmp[4182]*kernel[6]+tmp[4183]*kernel[7]+tmp[4184]*kernel[8];
				ans[4084]<=tmp[3983]*kernel[0]+tmp[3984]*kernel[1]+tmp[3985]*kernel[2]+tmp[4083]*kernel[3]+tmp[4084]*kernel[4]+tmp[4085]*kernel[5]+tmp[4183]*kernel[6]+tmp[4184]*kernel[7]+tmp[4185]*kernel[8];
				ans[4085]<=tmp[3984]*kernel[0]+tmp[3985]*kernel[1]+tmp[3986]*kernel[2]+tmp[4084]*kernel[3]+tmp[4085]*kernel[4]+tmp[4086]*kernel[5]+tmp[4184]*kernel[6]+tmp[4185]*kernel[7]+tmp[4186]*kernel[8];
				ans[4086]<=tmp[3985]*kernel[0]+tmp[3986]*kernel[1]+tmp[3987]*kernel[2]+tmp[4085]*kernel[3]+tmp[4086]*kernel[4]+tmp[4087]*kernel[5]+tmp[4185]*kernel[6]+tmp[4186]*kernel[7]+tmp[4187]*kernel[8];
				ans[4087]<=tmp[3986]*kernel[0]+tmp[3987]*kernel[1]+tmp[3988]*kernel[2]+tmp[4086]*kernel[3]+tmp[4087]*kernel[4]+tmp[4088]*kernel[5]+tmp[4186]*kernel[6]+tmp[4187]*kernel[7]+tmp[4188]*kernel[8];
				ans[4088]<=tmp[3987]*kernel[0]+tmp[3988]*kernel[1]+tmp[3989]*kernel[2]+tmp[4087]*kernel[3]+tmp[4088]*kernel[4]+tmp[4089]*kernel[5]+tmp[4187]*kernel[6]+tmp[4188]*kernel[7]+tmp[4189]*kernel[8];
				ans[4089]<=tmp[3988]*kernel[0]+tmp[3989]*kernel[1]+tmp[3990]*kernel[2]+tmp[4088]*kernel[3]+tmp[4089]*kernel[4]+tmp[4090]*kernel[5]+tmp[4188]*kernel[6]+tmp[4189]*kernel[7]+tmp[4190]*kernel[8];
				ans[4090]<=tmp[3989]*kernel[0]+tmp[3990]*kernel[1]+tmp[3991]*kernel[2]+tmp[4089]*kernel[3]+tmp[4090]*kernel[4]+tmp[4091]*kernel[5]+tmp[4189]*kernel[6]+tmp[4190]*kernel[7]+tmp[4191]*kernel[8];
				ans[4091]<=tmp[3990]*kernel[0]+tmp[3991]*kernel[1]+tmp[3992]*kernel[2]+tmp[4090]*kernel[3]+tmp[4091]*kernel[4]+tmp[4092]*kernel[5]+tmp[4190]*kernel[6]+tmp[4191]*kernel[7]+tmp[4192]*kernel[8];
				ans[4092]<=tmp[3991]*kernel[0]+tmp[3992]*kernel[1]+tmp[3993]*kernel[2]+tmp[4091]*kernel[3]+tmp[4092]*kernel[4]+tmp[4093]*kernel[5]+tmp[4191]*kernel[6]+tmp[4192]*kernel[7]+tmp[4193]*kernel[8];
				ans[4093]<=tmp[3992]*kernel[0]+tmp[3993]*kernel[1]+tmp[3994]*kernel[2]+tmp[4092]*kernel[3]+tmp[4093]*kernel[4]+tmp[4094]*kernel[5]+tmp[4192]*kernel[6]+tmp[4193]*kernel[7]+tmp[4194]*kernel[8];
				ans[4094]<=tmp[3993]*kernel[0]+tmp[3994]*kernel[1]+tmp[3995]*kernel[2]+tmp[4093]*kernel[3]+tmp[4094]*kernel[4]+tmp[4095]*kernel[5]+tmp[4193]*kernel[6]+tmp[4194]*kernel[7]+tmp[4195]*kernel[8];
				ans[4095]<=tmp[3994]*kernel[0]+tmp[3995]*kernel[1]+tmp[3996]*kernel[2]+tmp[4094]*kernel[3]+tmp[4095]*kernel[4]+tmp[4096]*kernel[5]+tmp[4194]*kernel[6]+tmp[4195]*kernel[7]+tmp[4196]*kernel[8];
				ans[4096]<=tmp[3995]*kernel[0]+tmp[3996]*kernel[1]+tmp[3997]*kernel[2]+tmp[4095]*kernel[3]+tmp[4096]*kernel[4]+tmp[4097]*kernel[5]+tmp[4195]*kernel[6]+tmp[4196]*kernel[7]+tmp[4197]*kernel[8];
				ans[4097]<=tmp[3996]*kernel[0]+tmp[3997]*kernel[1]+tmp[3998]*kernel[2]+tmp[4096]*kernel[3]+tmp[4097]*kernel[4]+tmp[4098]*kernel[5]+tmp[4196]*kernel[6]+tmp[4197]*kernel[7]+tmp[4198]*kernel[8];
				ans[4098]<=tmp[3997]*kernel[0]+tmp[3998]*kernel[1]+tmp[3999]*kernel[2]+tmp[4097]*kernel[3]+tmp[4098]*kernel[4]+tmp[4099]*kernel[5]+tmp[4197]*kernel[6]+tmp[4198]*kernel[7]+tmp[4199]*kernel[8];
				ans[4099]<=tmp[3998]*kernel[0]+tmp[3999]*kernel[1]+tmp[4098]*kernel[3]+tmp[4099]*kernel[4]+tmp[4198]*kernel[6]+tmp[4199]*kernel[7];
				ans[4100]<=tmp[4000]*kernel[1]+tmp[4001]*kernel[2]+tmp[4100]*kernel[4]+tmp[4101]*kernel[5]+tmp[4200]*kernel[7]+tmp[4201]*kernel[8];
				ans[4101]<=tmp[4000]*kernel[0]+tmp[4001]*kernel[1]+tmp[4002]*kernel[2]+tmp[4100]*kernel[3]+tmp[4101]*kernel[4]+tmp[4102]*kernel[5]+tmp[4200]*kernel[6]+tmp[4201]*kernel[7]+tmp[4202]*kernel[8];
				ans[4102]<=tmp[4001]*kernel[0]+tmp[4002]*kernel[1]+tmp[4003]*kernel[2]+tmp[4101]*kernel[3]+tmp[4102]*kernel[4]+tmp[4103]*kernel[5]+tmp[4201]*kernel[6]+tmp[4202]*kernel[7]+tmp[4203]*kernel[8];
				ans[4103]<=tmp[4002]*kernel[0]+tmp[4003]*kernel[1]+tmp[4004]*kernel[2]+tmp[4102]*kernel[3]+tmp[4103]*kernel[4]+tmp[4104]*kernel[5]+tmp[4202]*kernel[6]+tmp[4203]*kernel[7]+tmp[4204]*kernel[8];
				ans[4104]<=tmp[4003]*kernel[0]+tmp[4004]*kernel[1]+tmp[4005]*kernel[2]+tmp[4103]*kernel[3]+tmp[4104]*kernel[4]+tmp[4105]*kernel[5]+tmp[4203]*kernel[6]+tmp[4204]*kernel[7]+tmp[4205]*kernel[8];
				ans[4105]<=tmp[4004]*kernel[0]+tmp[4005]*kernel[1]+tmp[4006]*kernel[2]+tmp[4104]*kernel[3]+tmp[4105]*kernel[4]+tmp[4106]*kernel[5]+tmp[4204]*kernel[6]+tmp[4205]*kernel[7]+tmp[4206]*kernel[8];
				ans[4106]<=tmp[4005]*kernel[0]+tmp[4006]*kernel[1]+tmp[4007]*kernel[2]+tmp[4105]*kernel[3]+tmp[4106]*kernel[4]+tmp[4107]*kernel[5]+tmp[4205]*kernel[6]+tmp[4206]*kernel[7]+tmp[4207]*kernel[8];
				ans[4107]<=tmp[4006]*kernel[0]+tmp[4007]*kernel[1]+tmp[4008]*kernel[2]+tmp[4106]*kernel[3]+tmp[4107]*kernel[4]+tmp[4108]*kernel[5]+tmp[4206]*kernel[6]+tmp[4207]*kernel[7]+tmp[4208]*kernel[8];
				ans[4108]<=tmp[4007]*kernel[0]+tmp[4008]*kernel[1]+tmp[4009]*kernel[2]+tmp[4107]*kernel[3]+tmp[4108]*kernel[4]+tmp[4109]*kernel[5]+tmp[4207]*kernel[6]+tmp[4208]*kernel[7]+tmp[4209]*kernel[8];
				ans[4109]<=tmp[4008]*kernel[0]+tmp[4009]*kernel[1]+tmp[4010]*kernel[2]+tmp[4108]*kernel[3]+tmp[4109]*kernel[4]+tmp[4110]*kernel[5]+tmp[4208]*kernel[6]+tmp[4209]*kernel[7]+tmp[4210]*kernel[8];
				ans[4110]<=tmp[4009]*kernel[0]+tmp[4010]*kernel[1]+tmp[4011]*kernel[2]+tmp[4109]*kernel[3]+tmp[4110]*kernel[4]+tmp[4111]*kernel[5]+tmp[4209]*kernel[6]+tmp[4210]*kernel[7]+tmp[4211]*kernel[8];
				ans[4111]<=tmp[4010]*kernel[0]+tmp[4011]*kernel[1]+tmp[4012]*kernel[2]+tmp[4110]*kernel[3]+tmp[4111]*kernel[4]+tmp[4112]*kernel[5]+tmp[4210]*kernel[6]+tmp[4211]*kernel[7]+tmp[4212]*kernel[8];
				ans[4112]<=tmp[4011]*kernel[0]+tmp[4012]*kernel[1]+tmp[4013]*kernel[2]+tmp[4111]*kernel[3]+tmp[4112]*kernel[4]+tmp[4113]*kernel[5]+tmp[4211]*kernel[6]+tmp[4212]*kernel[7]+tmp[4213]*kernel[8];
				ans[4113]<=tmp[4012]*kernel[0]+tmp[4013]*kernel[1]+tmp[4014]*kernel[2]+tmp[4112]*kernel[3]+tmp[4113]*kernel[4]+tmp[4114]*kernel[5]+tmp[4212]*kernel[6]+tmp[4213]*kernel[7]+tmp[4214]*kernel[8];
				ans[4114]<=tmp[4013]*kernel[0]+tmp[4014]*kernel[1]+tmp[4015]*kernel[2]+tmp[4113]*kernel[3]+tmp[4114]*kernel[4]+tmp[4115]*kernel[5]+tmp[4213]*kernel[6]+tmp[4214]*kernel[7]+tmp[4215]*kernel[8];
				ans[4115]<=tmp[4014]*kernel[0]+tmp[4015]*kernel[1]+tmp[4016]*kernel[2]+tmp[4114]*kernel[3]+tmp[4115]*kernel[4]+tmp[4116]*kernel[5]+tmp[4214]*kernel[6]+tmp[4215]*kernel[7]+tmp[4216]*kernel[8];
				ans[4116]<=tmp[4015]*kernel[0]+tmp[4016]*kernel[1]+tmp[4017]*kernel[2]+tmp[4115]*kernel[3]+tmp[4116]*kernel[4]+tmp[4117]*kernel[5]+tmp[4215]*kernel[6]+tmp[4216]*kernel[7]+tmp[4217]*kernel[8];
				ans[4117]<=tmp[4016]*kernel[0]+tmp[4017]*kernel[1]+tmp[4018]*kernel[2]+tmp[4116]*kernel[3]+tmp[4117]*kernel[4]+tmp[4118]*kernel[5]+tmp[4216]*kernel[6]+tmp[4217]*kernel[7]+tmp[4218]*kernel[8];
				ans[4118]<=tmp[4017]*kernel[0]+tmp[4018]*kernel[1]+tmp[4019]*kernel[2]+tmp[4117]*kernel[3]+tmp[4118]*kernel[4]+tmp[4119]*kernel[5]+tmp[4217]*kernel[6]+tmp[4218]*kernel[7]+tmp[4219]*kernel[8];
				ans[4119]<=tmp[4018]*kernel[0]+tmp[4019]*kernel[1]+tmp[4020]*kernel[2]+tmp[4118]*kernel[3]+tmp[4119]*kernel[4]+tmp[4120]*kernel[5]+tmp[4218]*kernel[6]+tmp[4219]*kernel[7]+tmp[4220]*kernel[8];
				ans[4120]<=tmp[4019]*kernel[0]+tmp[4020]*kernel[1]+tmp[4021]*kernel[2]+tmp[4119]*kernel[3]+tmp[4120]*kernel[4]+tmp[4121]*kernel[5]+tmp[4219]*kernel[6]+tmp[4220]*kernel[7]+tmp[4221]*kernel[8];
				ans[4121]<=tmp[4020]*kernel[0]+tmp[4021]*kernel[1]+tmp[4022]*kernel[2]+tmp[4120]*kernel[3]+tmp[4121]*kernel[4]+tmp[4122]*kernel[5]+tmp[4220]*kernel[6]+tmp[4221]*kernel[7]+tmp[4222]*kernel[8];
				ans[4122]<=tmp[4021]*kernel[0]+tmp[4022]*kernel[1]+tmp[4023]*kernel[2]+tmp[4121]*kernel[3]+tmp[4122]*kernel[4]+tmp[4123]*kernel[5]+tmp[4221]*kernel[6]+tmp[4222]*kernel[7]+tmp[4223]*kernel[8];
				ans[4123]<=tmp[4022]*kernel[0]+tmp[4023]*kernel[1]+tmp[4024]*kernel[2]+tmp[4122]*kernel[3]+tmp[4123]*kernel[4]+tmp[4124]*kernel[5]+tmp[4222]*kernel[6]+tmp[4223]*kernel[7]+tmp[4224]*kernel[8];
				ans[4124]<=tmp[4023]*kernel[0]+tmp[4024]*kernel[1]+tmp[4025]*kernel[2]+tmp[4123]*kernel[3]+tmp[4124]*kernel[4]+tmp[4125]*kernel[5]+tmp[4223]*kernel[6]+tmp[4224]*kernel[7]+tmp[4225]*kernel[8];
				ans[4125]<=tmp[4024]*kernel[0]+tmp[4025]*kernel[1]+tmp[4026]*kernel[2]+tmp[4124]*kernel[3]+tmp[4125]*kernel[4]+tmp[4126]*kernel[5]+tmp[4224]*kernel[6]+tmp[4225]*kernel[7]+tmp[4226]*kernel[8];
				ans[4126]<=tmp[4025]*kernel[0]+tmp[4026]*kernel[1]+tmp[4027]*kernel[2]+tmp[4125]*kernel[3]+tmp[4126]*kernel[4]+tmp[4127]*kernel[5]+tmp[4225]*kernel[6]+tmp[4226]*kernel[7]+tmp[4227]*kernel[8];
				ans[4127]<=tmp[4026]*kernel[0]+tmp[4027]*kernel[1]+tmp[4028]*kernel[2]+tmp[4126]*kernel[3]+tmp[4127]*kernel[4]+tmp[4128]*kernel[5]+tmp[4226]*kernel[6]+tmp[4227]*kernel[7]+tmp[4228]*kernel[8];
				ans[4128]<=tmp[4027]*kernel[0]+tmp[4028]*kernel[1]+tmp[4029]*kernel[2]+tmp[4127]*kernel[3]+tmp[4128]*kernel[4]+tmp[4129]*kernel[5]+tmp[4227]*kernel[6]+tmp[4228]*kernel[7]+tmp[4229]*kernel[8];
				ans[4129]<=tmp[4028]*kernel[0]+tmp[4029]*kernel[1]+tmp[4030]*kernel[2]+tmp[4128]*kernel[3]+tmp[4129]*kernel[4]+tmp[4130]*kernel[5]+tmp[4228]*kernel[6]+tmp[4229]*kernel[7]+tmp[4230]*kernel[8];
				ans[4130]<=tmp[4029]*kernel[0]+tmp[4030]*kernel[1]+tmp[4031]*kernel[2]+tmp[4129]*kernel[3]+tmp[4130]*kernel[4]+tmp[4131]*kernel[5]+tmp[4229]*kernel[6]+tmp[4230]*kernel[7]+tmp[4231]*kernel[8];
				ans[4131]<=tmp[4030]*kernel[0]+tmp[4031]*kernel[1]+tmp[4032]*kernel[2]+tmp[4130]*kernel[3]+tmp[4131]*kernel[4]+tmp[4132]*kernel[5]+tmp[4230]*kernel[6]+tmp[4231]*kernel[7]+tmp[4232]*kernel[8];
				ans[4132]<=tmp[4031]*kernel[0]+tmp[4032]*kernel[1]+tmp[4033]*kernel[2]+tmp[4131]*kernel[3]+tmp[4132]*kernel[4]+tmp[4133]*kernel[5]+tmp[4231]*kernel[6]+tmp[4232]*kernel[7]+tmp[4233]*kernel[8];
				ans[4133]<=tmp[4032]*kernel[0]+tmp[4033]*kernel[1]+tmp[4034]*kernel[2]+tmp[4132]*kernel[3]+tmp[4133]*kernel[4]+tmp[4134]*kernel[5]+tmp[4232]*kernel[6]+tmp[4233]*kernel[7]+tmp[4234]*kernel[8];
				ans[4134]<=tmp[4033]*kernel[0]+tmp[4034]*kernel[1]+tmp[4035]*kernel[2]+tmp[4133]*kernel[3]+tmp[4134]*kernel[4]+tmp[4135]*kernel[5]+tmp[4233]*kernel[6]+tmp[4234]*kernel[7]+tmp[4235]*kernel[8];
				ans[4135]<=tmp[4034]*kernel[0]+tmp[4035]*kernel[1]+tmp[4036]*kernel[2]+tmp[4134]*kernel[3]+tmp[4135]*kernel[4]+tmp[4136]*kernel[5]+tmp[4234]*kernel[6]+tmp[4235]*kernel[7]+tmp[4236]*kernel[8];
				ans[4136]<=tmp[4035]*kernel[0]+tmp[4036]*kernel[1]+tmp[4037]*kernel[2]+tmp[4135]*kernel[3]+tmp[4136]*kernel[4]+tmp[4137]*kernel[5]+tmp[4235]*kernel[6]+tmp[4236]*kernel[7]+tmp[4237]*kernel[8];
				ans[4137]<=tmp[4036]*kernel[0]+tmp[4037]*kernel[1]+tmp[4038]*kernel[2]+tmp[4136]*kernel[3]+tmp[4137]*kernel[4]+tmp[4138]*kernel[5]+tmp[4236]*kernel[6]+tmp[4237]*kernel[7]+tmp[4238]*kernel[8];
				ans[4138]<=tmp[4037]*kernel[0]+tmp[4038]*kernel[1]+tmp[4039]*kernel[2]+tmp[4137]*kernel[3]+tmp[4138]*kernel[4]+tmp[4139]*kernel[5]+tmp[4237]*kernel[6]+tmp[4238]*kernel[7]+tmp[4239]*kernel[8];
				ans[4139]<=tmp[4038]*kernel[0]+tmp[4039]*kernel[1]+tmp[4040]*kernel[2]+tmp[4138]*kernel[3]+tmp[4139]*kernel[4]+tmp[4140]*kernel[5]+tmp[4238]*kernel[6]+tmp[4239]*kernel[7]+tmp[4240]*kernel[8];
				ans[4140]<=tmp[4039]*kernel[0]+tmp[4040]*kernel[1]+tmp[4041]*kernel[2]+tmp[4139]*kernel[3]+tmp[4140]*kernel[4]+tmp[4141]*kernel[5]+tmp[4239]*kernel[6]+tmp[4240]*kernel[7]+tmp[4241]*kernel[8];
				ans[4141]<=tmp[4040]*kernel[0]+tmp[4041]*kernel[1]+tmp[4042]*kernel[2]+tmp[4140]*kernel[3]+tmp[4141]*kernel[4]+tmp[4142]*kernel[5]+tmp[4240]*kernel[6]+tmp[4241]*kernel[7]+tmp[4242]*kernel[8];
				ans[4142]<=tmp[4041]*kernel[0]+tmp[4042]*kernel[1]+tmp[4043]*kernel[2]+tmp[4141]*kernel[3]+tmp[4142]*kernel[4]+tmp[4143]*kernel[5]+tmp[4241]*kernel[6]+tmp[4242]*kernel[7]+tmp[4243]*kernel[8];
				ans[4143]<=tmp[4042]*kernel[0]+tmp[4043]*kernel[1]+tmp[4044]*kernel[2]+tmp[4142]*kernel[3]+tmp[4143]*kernel[4]+tmp[4144]*kernel[5]+tmp[4242]*kernel[6]+tmp[4243]*kernel[7]+tmp[4244]*kernel[8];
				ans[4144]<=tmp[4043]*kernel[0]+tmp[4044]*kernel[1]+tmp[4045]*kernel[2]+tmp[4143]*kernel[3]+tmp[4144]*kernel[4]+tmp[4145]*kernel[5]+tmp[4243]*kernel[6]+tmp[4244]*kernel[7]+tmp[4245]*kernel[8];
				ans[4145]<=tmp[4044]*kernel[0]+tmp[4045]*kernel[1]+tmp[4046]*kernel[2]+tmp[4144]*kernel[3]+tmp[4145]*kernel[4]+tmp[4146]*kernel[5]+tmp[4244]*kernel[6]+tmp[4245]*kernel[7]+tmp[4246]*kernel[8];
				ans[4146]<=tmp[4045]*kernel[0]+tmp[4046]*kernel[1]+tmp[4047]*kernel[2]+tmp[4145]*kernel[3]+tmp[4146]*kernel[4]+tmp[4147]*kernel[5]+tmp[4245]*kernel[6]+tmp[4246]*kernel[7]+tmp[4247]*kernel[8];
				ans[4147]<=tmp[4046]*kernel[0]+tmp[4047]*kernel[1]+tmp[4048]*kernel[2]+tmp[4146]*kernel[3]+tmp[4147]*kernel[4]+tmp[4148]*kernel[5]+tmp[4246]*kernel[6]+tmp[4247]*kernel[7]+tmp[4248]*kernel[8];
				ans[4148]<=tmp[4047]*kernel[0]+tmp[4048]*kernel[1]+tmp[4049]*kernel[2]+tmp[4147]*kernel[3]+tmp[4148]*kernel[4]+tmp[4149]*kernel[5]+tmp[4247]*kernel[6]+tmp[4248]*kernel[7]+tmp[4249]*kernel[8];
				ans[4149]<=tmp[4048]*kernel[0]+tmp[4049]*kernel[1]+tmp[4050]*kernel[2]+tmp[4148]*kernel[3]+tmp[4149]*kernel[4]+tmp[4150]*kernel[5]+tmp[4248]*kernel[6]+tmp[4249]*kernel[7]+tmp[4250]*kernel[8];
				ans[4150]<=tmp[4049]*kernel[0]+tmp[4050]*kernel[1]+tmp[4051]*kernel[2]+tmp[4149]*kernel[3]+tmp[4150]*kernel[4]+tmp[4151]*kernel[5]+tmp[4249]*kernel[6]+tmp[4250]*kernel[7]+tmp[4251]*kernel[8];
				ans[4151]<=tmp[4050]*kernel[0]+tmp[4051]*kernel[1]+tmp[4052]*kernel[2]+tmp[4150]*kernel[3]+tmp[4151]*kernel[4]+tmp[4152]*kernel[5]+tmp[4250]*kernel[6]+tmp[4251]*kernel[7]+tmp[4252]*kernel[8];
				ans[4152]<=tmp[4051]*kernel[0]+tmp[4052]*kernel[1]+tmp[4053]*kernel[2]+tmp[4151]*kernel[3]+tmp[4152]*kernel[4]+tmp[4153]*kernel[5]+tmp[4251]*kernel[6]+tmp[4252]*kernel[7]+tmp[4253]*kernel[8];
				ans[4153]<=tmp[4052]*kernel[0]+tmp[4053]*kernel[1]+tmp[4054]*kernel[2]+tmp[4152]*kernel[3]+tmp[4153]*kernel[4]+tmp[4154]*kernel[5]+tmp[4252]*kernel[6]+tmp[4253]*kernel[7]+tmp[4254]*kernel[8];
				ans[4154]<=tmp[4053]*kernel[0]+tmp[4054]*kernel[1]+tmp[4055]*kernel[2]+tmp[4153]*kernel[3]+tmp[4154]*kernel[4]+tmp[4155]*kernel[5]+tmp[4253]*kernel[6]+tmp[4254]*kernel[7]+tmp[4255]*kernel[8];
				ans[4155]<=tmp[4054]*kernel[0]+tmp[4055]*kernel[1]+tmp[4056]*kernel[2]+tmp[4154]*kernel[3]+tmp[4155]*kernel[4]+tmp[4156]*kernel[5]+tmp[4254]*kernel[6]+tmp[4255]*kernel[7]+tmp[4256]*kernel[8];
				ans[4156]<=tmp[4055]*kernel[0]+tmp[4056]*kernel[1]+tmp[4057]*kernel[2]+tmp[4155]*kernel[3]+tmp[4156]*kernel[4]+tmp[4157]*kernel[5]+tmp[4255]*kernel[6]+tmp[4256]*kernel[7]+tmp[4257]*kernel[8];
				ans[4157]<=tmp[4056]*kernel[0]+tmp[4057]*kernel[1]+tmp[4058]*kernel[2]+tmp[4156]*kernel[3]+tmp[4157]*kernel[4]+tmp[4158]*kernel[5]+tmp[4256]*kernel[6]+tmp[4257]*kernel[7]+tmp[4258]*kernel[8];
				ans[4158]<=tmp[4057]*kernel[0]+tmp[4058]*kernel[1]+tmp[4059]*kernel[2]+tmp[4157]*kernel[3]+tmp[4158]*kernel[4]+tmp[4159]*kernel[5]+tmp[4257]*kernel[6]+tmp[4258]*kernel[7]+tmp[4259]*kernel[8];
				ans[4159]<=tmp[4058]*kernel[0]+tmp[4059]*kernel[1]+tmp[4060]*kernel[2]+tmp[4158]*kernel[3]+tmp[4159]*kernel[4]+tmp[4160]*kernel[5]+tmp[4258]*kernel[6]+tmp[4259]*kernel[7]+tmp[4260]*kernel[8];
				ans[4160]<=tmp[4059]*kernel[0]+tmp[4060]*kernel[1]+tmp[4061]*kernel[2]+tmp[4159]*kernel[3]+tmp[4160]*kernel[4]+tmp[4161]*kernel[5]+tmp[4259]*kernel[6]+tmp[4260]*kernel[7]+tmp[4261]*kernel[8];
				ans[4161]<=tmp[4060]*kernel[0]+tmp[4061]*kernel[1]+tmp[4062]*kernel[2]+tmp[4160]*kernel[3]+tmp[4161]*kernel[4]+tmp[4162]*kernel[5]+tmp[4260]*kernel[6]+tmp[4261]*kernel[7]+tmp[4262]*kernel[8];
				ans[4162]<=tmp[4061]*kernel[0]+tmp[4062]*kernel[1]+tmp[4063]*kernel[2]+tmp[4161]*kernel[3]+tmp[4162]*kernel[4]+tmp[4163]*kernel[5]+tmp[4261]*kernel[6]+tmp[4262]*kernel[7]+tmp[4263]*kernel[8];
				ans[4163]<=tmp[4062]*kernel[0]+tmp[4063]*kernel[1]+tmp[4064]*kernel[2]+tmp[4162]*kernel[3]+tmp[4163]*kernel[4]+tmp[4164]*kernel[5]+tmp[4262]*kernel[6]+tmp[4263]*kernel[7]+tmp[4264]*kernel[8];
				ans[4164]<=tmp[4063]*kernel[0]+tmp[4064]*kernel[1]+tmp[4065]*kernel[2]+tmp[4163]*kernel[3]+tmp[4164]*kernel[4]+tmp[4165]*kernel[5]+tmp[4263]*kernel[6]+tmp[4264]*kernel[7]+tmp[4265]*kernel[8];
				ans[4165]<=tmp[4064]*kernel[0]+tmp[4065]*kernel[1]+tmp[4066]*kernel[2]+tmp[4164]*kernel[3]+tmp[4165]*kernel[4]+tmp[4166]*kernel[5]+tmp[4264]*kernel[6]+tmp[4265]*kernel[7]+tmp[4266]*kernel[8];
				ans[4166]<=tmp[4065]*kernel[0]+tmp[4066]*kernel[1]+tmp[4067]*kernel[2]+tmp[4165]*kernel[3]+tmp[4166]*kernel[4]+tmp[4167]*kernel[5]+tmp[4265]*kernel[6]+tmp[4266]*kernel[7]+tmp[4267]*kernel[8];
				ans[4167]<=tmp[4066]*kernel[0]+tmp[4067]*kernel[1]+tmp[4068]*kernel[2]+tmp[4166]*kernel[3]+tmp[4167]*kernel[4]+tmp[4168]*kernel[5]+tmp[4266]*kernel[6]+tmp[4267]*kernel[7]+tmp[4268]*kernel[8];
				ans[4168]<=tmp[4067]*kernel[0]+tmp[4068]*kernel[1]+tmp[4069]*kernel[2]+tmp[4167]*kernel[3]+tmp[4168]*kernel[4]+tmp[4169]*kernel[5]+tmp[4267]*kernel[6]+tmp[4268]*kernel[7]+tmp[4269]*kernel[8];
				ans[4169]<=tmp[4068]*kernel[0]+tmp[4069]*kernel[1]+tmp[4070]*kernel[2]+tmp[4168]*kernel[3]+tmp[4169]*kernel[4]+tmp[4170]*kernel[5]+tmp[4268]*kernel[6]+tmp[4269]*kernel[7]+tmp[4270]*kernel[8];
				ans[4170]<=tmp[4069]*kernel[0]+tmp[4070]*kernel[1]+tmp[4071]*kernel[2]+tmp[4169]*kernel[3]+tmp[4170]*kernel[4]+tmp[4171]*kernel[5]+tmp[4269]*kernel[6]+tmp[4270]*kernel[7]+tmp[4271]*kernel[8];
				ans[4171]<=tmp[4070]*kernel[0]+tmp[4071]*kernel[1]+tmp[4072]*kernel[2]+tmp[4170]*kernel[3]+tmp[4171]*kernel[4]+tmp[4172]*kernel[5]+tmp[4270]*kernel[6]+tmp[4271]*kernel[7]+tmp[4272]*kernel[8];
				ans[4172]<=tmp[4071]*kernel[0]+tmp[4072]*kernel[1]+tmp[4073]*kernel[2]+tmp[4171]*kernel[3]+tmp[4172]*kernel[4]+tmp[4173]*kernel[5]+tmp[4271]*kernel[6]+tmp[4272]*kernel[7]+tmp[4273]*kernel[8];
				ans[4173]<=tmp[4072]*kernel[0]+tmp[4073]*kernel[1]+tmp[4074]*kernel[2]+tmp[4172]*kernel[3]+tmp[4173]*kernel[4]+tmp[4174]*kernel[5]+tmp[4272]*kernel[6]+tmp[4273]*kernel[7]+tmp[4274]*kernel[8];
				ans[4174]<=tmp[4073]*kernel[0]+tmp[4074]*kernel[1]+tmp[4075]*kernel[2]+tmp[4173]*kernel[3]+tmp[4174]*kernel[4]+tmp[4175]*kernel[5]+tmp[4273]*kernel[6]+tmp[4274]*kernel[7]+tmp[4275]*kernel[8];
				ans[4175]<=tmp[4074]*kernel[0]+tmp[4075]*kernel[1]+tmp[4076]*kernel[2]+tmp[4174]*kernel[3]+tmp[4175]*kernel[4]+tmp[4176]*kernel[5]+tmp[4274]*kernel[6]+tmp[4275]*kernel[7]+tmp[4276]*kernel[8];
				ans[4176]<=tmp[4075]*kernel[0]+tmp[4076]*kernel[1]+tmp[4077]*kernel[2]+tmp[4175]*kernel[3]+tmp[4176]*kernel[4]+tmp[4177]*kernel[5]+tmp[4275]*kernel[6]+tmp[4276]*kernel[7]+tmp[4277]*kernel[8];
				ans[4177]<=tmp[4076]*kernel[0]+tmp[4077]*kernel[1]+tmp[4078]*kernel[2]+tmp[4176]*kernel[3]+tmp[4177]*kernel[4]+tmp[4178]*kernel[5]+tmp[4276]*kernel[6]+tmp[4277]*kernel[7]+tmp[4278]*kernel[8];
				ans[4178]<=tmp[4077]*kernel[0]+tmp[4078]*kernel[1]+tmp[4079]*kernel[2]+tmp[4177]*kernel[3]+tmp[4178]*kernel[4]+tmp[4179]*kernel[5]+tmp[4277]*kernel[6]+tmp[4278]*kernel[7]+tmp[4279]*kernel[8];
				ans[4179]<=tmp[4078]*kernel[0]+tmp[4079]*kernel[1]+tmp[4080]*kernel[2]+tmp[4178]*kernel[3]+tmp[4179]*kernel[4]+tmp[4180]*kernel[5]+tmp[4278]*kernel[6]+tmp[4279]*kernel[7]+tmp[4280]*kernel[8];
				ans[4180]<=tmp[4079]*kernel[0]+tmp[4080]*kernel[1]+tmp[4081]*kernel[2]+tmp[4179]*kernel[3]+tmp[4180]*kernel[4]+tmp[4181]*kernel[5]+tmp[4279]*kernel[6]+tmp[4280]*kernel[7]+tmp[4281]*kernel[8];
				ans[4181]<=tmp[4080]*kernel[0]+tmp[4081]*kernel[1]+tmp[4082]*kernel[2]+tmp[4180]*kernel[3]+tmp[4181]*kernel[4]+tmp[4182]*kernel[5]+tmp[4280]*kernel[6]+tmp[4281]*kernel[7]+tmp[4282]*kernel[8];
				ans[4182]<=tmp[4081]*kernel[0]+tmp[4082]*kernel[1]+tmp[4083]*kernel[2]+tmp[4181]*kernel[3]+tmp[4182]*kernel[4]+tmp[4183]*kernel[5]+tmp[4281]*kernel[6]+tmp[4282]*kernel[7]+tmp[4283]*kernel[8];
				ans[4183]<=tmp[4082]*kernel[0]+tmp[4083]*kernel[1]+tmp[4084]*kernel[2]+tmp[4182]*kernel[3]+tmp[4183]*kernel[4]+tmp[4184]*kernel[5]+tmp[4282]*kernel[6]+tmp[4283]*kernel[7]+tmp[4284]*kernel[8];
				ans[4184]<=tmp[4083]*kernel[0]+tmp[4084]*kernel[1]+tmp[4085]*kernel[2]+tmp[4183]*kernel[3]+tmp[4184]*kernel[4]+tmp[4185]*kernel[5]+tmp[4283]*kernel[6]+tmp[4284]*kernel[7]+tmp[4285]*kernel[8];
				ans[4185]<=tmp[4084]*kernel[0]+tmp[4085]*kernel[1]+tmp[4086]*kernel[2]+tmp[4184]*kernel[3]+tmp[4185]*kernel[4]+tmp[4186]*kernel[5]+tmp[4284]*kernel[6]+tmp[4285]*kernel[7]+tmp[4286]*kernel[8];
				ans[4186]<=tmp[4085]*kernel[0]+tmp[4086]*kernel[1]+tmp[4087]*kernel[2]+tmp[4185]*kernel[3]+tmp[4186]*kernel[4]+tmp[4187]*kernel[5]+tmp[4285]*kernel[6]+tmp[4286]*kernel[7]+tmp[4287]*kernel[8];
				ans[4187]<=tmp[4086]*kernel[0]+tmp[4087]*kernel[1]+tmp[4088]*kernel[2]+tmp[4186]*kernel[3]+tmp[4187]*kernel[4]+tmp[4188]*kernel[5]+tmp[4286]*kernel[6]+tmp[4287]*kernel[7]+tmp[4288]*kernel[8];
				ans[4188]<=tmp[4087]*kernel[0]+tmp[4088]*kernel[1]+tmp[4089]*kernel[2]+tmp[4187]*kernel[3]+tmp[4188]*kernel[4]+tmp[4189]*kernel[5]+tmp[4287]*kernel[6]+tmp[4288]*kernel[7]+tmp[4289]*kernel[8];
				ans[4189]<=tmp[4088]*kernel[0]+tmp[4089]*kernel[1]+tmp[4090]*kernel[2]+tmp[4188]*kernel[3]+tmp[4189]*kernel[4]+tmp[4190]*kernel[5]+tmp[4288]*kernel[6]+tmp[4289]*kernel[7]+tmp[4290]*kernel[8];
				ans[4190]<=tmp[4089]*kernel[0]+tmp[4090]*kernel[1]+tmp[4091]*kernel[2]+tmp[4189]*kernel[3]+tmp[4190]*kernel[4]+tmp[4191]*kernel[5]+tmp[4289]*kernel[6]+tmp[4290]*kernel[7]+tmp[4291]*kernel[8];
				ans[4191]<=tmp[4090]*kernel[0]+tmp[4091]*kernel[1]+tmp[4092]*kernel[2]+tmp[4190]*kernel[3]+tmp[4191]*kernel[4]+tmp[4192]*kernel[5]+tmp[4290]*kernel[6]+tmp[4291]*kernel[7]+tmp[4292]*kernel[8];
				ans[4192]<=tmp[4091]*kernel[0]+tmp[4092]*kernel[1]+tmp[4093]*kernel[2]+tmp[4191]*kernel[3]+tmp[4192]*kernel[4]+tmp[4193]*kernel[5]+tmp[4291]*kernel[6]+tmp[4292]*kernel[7]+tmp[4293]*kernel[8];
				ans[4193]<=tmp[4092]*kernel[0]+tmp[4093]*kernel[1]+tmp[4094]*kernel[2]+tmp[4192]*kernel[3]+tmp[4193]*kernel[4]+tmp[4194]*kernel[5]+tmp[4292]*kernel[6]+tmp[4293]*kernel[7]+tmp[4294]*kernel[8];
				ans[4194]<=tmp[4093]*kernel[0]+tmp[4094]*kernel[1]+tmp[4095]*kernel[2]+tmp[4193]*kernel[3]+tmp[4194]*kernel[4]+tmp[4195]*kernel[5]+tmp[4293]*kernel[6]+tmp[4294]*kernel[7]+tmp[4295]*kernel[8];
				ans[4195]<=tmp[4094]*kernel[0]+tmp[4095]*kernel[1]+tmp[4096]*kernel[2]+tmp[4194]*kernel[3]+tmp[4195]*kernel[4]+tmp[4196]*kernel[5]+tmp[4294]*kernel[6]+tmp[4295]*kernel[7]+tmp[4296]*kernel[8];
				ans[4196]<=tmp[4095]*kernel[0]+tmp[4096]*kernel[1]+tmp[4097]*kernel[2]+tmp[4195]*kernel[3]+tmp[4196]*kernel[4]+tmp[4197]*kernel[5]+tmp[4295]*kernel[6]+tmp[4296]*kernel[7]+tmp[4297]*kernel[8];
				ans[4197]<=tmp[4096]*kernel[0]+tmp[4097]*kernel[1]+tmp[4098]*kernel[2]+tmp[4196]*kernel[3]+tmp[4197]*kernel[4]+tmp[4198]*kernel[5]+tmp[4296]*kernel[6]+tmp[4297]*kernel[7]+tmp[4298]*kernel[8];
				ans[4198]<=tmp[4097]*kernel[0]+tmp[4098]*kernel[1]+tmp[4099]*kernel[2]+tmp[4197]*kernel[3]+tmp[4198]*kernel[4]+tmp[4199]*kernel[5]+tmp[4297]*kernel[6]+tmp[4298]*kernel[7]+tmp[4299]*kernel[8];
				ans[4199]<=tmp[4098]*kernel[0]+tmp[4099]*kernel[1]+tmp[4198]*kernel[3]+tmp[4199]*kernel[4]+tmp[4298]*kernel[6]+tmp[4299]*kernel[7];
				ans[4200]<=tmp[4100]*kernel[1]+tmp[4101]*kernel[2]+tmp[4200]*kernel[4]+tmp[4201]*kernel[5]+tmp[4300]*kernel[7]+tmp[4301]*kernel[8];
				ans[4201]<=tmp[4100]*kernel[0]+tmp[4101]*kernel[1]+tmp[4102]*kernel[2]+tmp[4200]*kernel[3]+tmp[4201]*kernel[4]+tmp[4202]*kernel[5]+tmp[4300]*kernel[6]+tmp[4301]*kernel[7]+tmp[4302]*kernel[8];
				ans[4202]<=tmp[4101]*kernel[0]+tmp[4102]*kernel[1]+tmp[4103]*kernel[2]+tmp[4201]*kernel[3]+tmp[4202]*kernel[4]+tmp[4203]*kernel[5]+tmp[4301]*kernel[6]+tmp[4302]*kernel[7]+tmp[4303]*kernel[8];
				ans[4203]<=tmp[4102]*kernel[0]+tmp[4103]*kernel[1]+tmp[4104]*kernel[2]+tmp[4202]*kernel[3]+tmp[4203]*kernel[4]+tmp[4204]*kernel[5]+tmp[4302]*kernel[6]+tmp[4303]*kernel[7]+tmp[4304]*kernel[8];
				ans[4204]<=tmp[4103]*kernel[0]+tmp[4104]*kernel[1]+tmp[4105]*kernel[2]+tmp[4203]*kernel[3]+tmp[4204]*kernel[4]+tmp[4205]*kernel[5]+tmp[4303]*kernel[6]+tmp[4304]*kernel[7]+tmp[4305]*kernel[8];
				ans[4205]<=tmp[4104]*kernel[0]+tmp[4105]*kernel[1]+tmp[4106]*kernel[2]+tmp[4204]*kernel[3]+tmp[4205]*kernel[4]+tmp[4206]*kernel[5]+tmp[4304]*kernel[6]+tmp[4305]*kernel[7]+tmp[4306]*kernel[8];
				ans[4206]<=tmp[4105]*kernel[0]+tmp[4106]*kernel[1]+tmp[4107]*kernel[2]+tmp[4205]*kernel[3]+tmp[4206]*kernel[4]+tmp[4207]*kernel[5]+tmp[4305]*kernel[6]+tmp[4306]*kernel[7]+tmp[4307]*kernel[8];
				ans[4207]<=tmp[4106]*kernel[0]+tmp[4107]*kernel[1]+tmp[4108]*kernel[2]+tmp[4206]*kernel[3]+tmp[4207]*kernel[4]+tmp[4208]*kernel[5]+tmp[4306]*kernel[6]+tmp[4307]*kernel[7]+tmp[4308]*kernel[8];
				ans[4208]<=tmp[4107]*kernel[0]+tmp[4108]*kernel[1]+tmp[4109]*kernel[2]+tmp[4207]*kernel[3]+tmp[4208]*kernel[4]+tmp[4209]*kernel[5]+tmp[4307]*kernel[6]+tmp[4308]*kernel[7]+tmp[4309]*kernel[8];
				ans[4209]<=tmp[4108]*kernel[0]+tmp[4109]*kernel[1]+tmp[4110]*kernel[2]+tmp[4208]*kernel[3]+tmp[4209]*kernel[4]+tmp[4210]*kernel[5]+tmp[4308]*kernel[6]+tmp[4309]*kernel[7]+tmp[4310]*kernel[8];
				ans[4210]<=tmp[4109]*kernel[0]+tmp[4110]*kernel[1]+tmp[4111]*kernel[2]+tmp[4209]*kernel[3]+tmp[4210]*kernel[4]+tmp[4211]*kernel[5]+tmp[4309]*kernel[6]+tmp[4310]*kernel[7]+tmp[4311]*kernel[8];
				ans[4211]<=tmp[4110]*kernel[0]+tmp[4111]*kernel[1]+tmp[4112]*kernel[2]+tmp[4210]*kernel[3]+tmp[4211]*kernel[4]+tmp[4212]*kernel[5]+tmp[4310]*kernel[6]+tmp[4311]*kernel[7]+tmp[4312]*kernel[8];
				ans[4212]<=tmp[4111]*kernel[0]+tmp[4112]*kernel[1]+tmp[4113]*kernel[2]+tmp[4211]*kernel[3]+tmp[4212]*kernel[4]+tmp[4213]*kernel[5]+tmp[4311]*kernel[6]+tmp[4312]*kernel[7]+tmp[4313]*kernel[8];
				ans[4213]<=tmp[4112]*kernel[0]+tmp[4113]*kernel[1]+tmp[4114]*kernel[2]+tmp[4212]*kernel[3]+tmp[4213]*kernel[4]+tmp[4214]*kernel[5]+tmp[4312]*kernel[6]+tmp[4313]*kernel[7]+tmp[4314]*kernel[8];
				ans[4214]<=tmp[4113]*kernel[0]+tmp[4114]*kernel[1]+tmp[4115]*kernel[2]+tmp[4213]*kernel[3]+tmp[4214]*kernel[4]+tmp[4215]*kernel[5]+tmp[4313]*kernel[6]+tmp[4314]*kernel[7]+tmp[4315]*kernel[8];
				ans[4215]<=tmp[4114]*kernel[0]+tmp[4115]*kernel[1]+tmp[4116]*kernel[2]+tmp[4214]*kernel[3]+tmp[4215]*kernel[4]+tmp[4216]*kernel[5]+tmp[4314]*kernel[6]+tmp[4315]*kernel[7]+tmp[4316]*kernel[8];
				ans[4216]<=tmp[4115]*kernel[0]+tmp[4116]*kernel[1]+tmp[4117]*kernel[2]+tmp[4215]*kernel[3]+tmp[4216]*kernel[4]+tmp[4217]*kernel[5]+tmp[4315]*kernel[6]+tmp[4316]*kernel[7]+tmp[4317]*kernel[8];
				ans[4217]<=tmp[4116]*kernel[0]+tmp[4117]*kernel[1]+tmp[4118]*kernel[2]+tmp[4216]*kernel[3]+tmp[4217]*kernel[4]+tmp[4218]*kernel[5]+tmp[4316]*kernel[6]+tmp[4317]*kernel[7]+tmp[4318]*kernel[8];
				ans[4218]<=tmp[4117]*kernel[0]+tmp[4118]*kernel[1]+tmp[4119]*kernel[2]+tmp[4217]*kernel[3]+tmp[4218]*kernel[4]+tmp[4219]*kernel[5]+tmp[4317]*kernel[6]+tmp[4318]*kernel[7]+tmp[4319]*kernel[8];
				ans[4219]<=tmp[4118]*kernel[0]+tmp[4119]*kernel[1]+tmp[4120]*kernel[2]+tmp[4218]*kernel[3]+tmp[4219]*kernel[4]+tmp[4220]*kernel[5]+tmp[4318]*kernel[6]+tmp[4319]*kernel[7]+tmp[4320]*kernel[8];
				ans[4220]<=tmp[4119]*kernel[0]+tmp[4120]*kernel[1]+tmp[4121]*kernel[2]+tmp[4219]*kernel[3]+tmp[4220]*kernel[4]+tmp[4221]*kernel[5]+tmp[4319]*kernel[6]+tmp[4320]*kernel[7]+tmp[4321]*kernel[8];
				ans[4221]<=tmp[4120]*kernel[0]+tmp[4121]*kernel[1]+tmp[4122]*kernel[2]+tmp[4220]*kernel[3]+tmp[4221]*kernel[4]+tmp[4222]*kernel[5]+tmp[4320]*kernel[6]+tmp[4321]*kernel[7]+tmp[4322]*kernel[8];
				ans[4222]<=tmp[4121]*kernel[0]+tmp[4122]*kernel[1]+tmp[4123]*kernel[2]+tmp[4221]*kernel[3]+tmp[4222]*kernel[4]+tmp[4223]*kernel[5]+tmp[4321]*kernel[6]+tmp[4322]*kernel[7]+tmp[4323]*kernel[8];
				ans[4223]<=tmp[4122]*kernel[0]+tmp[4123]*kernel[1]+tmp[4124]*kernel[2]+tmp[4222]*kernel[3]+tmp[4223]*kernel[4]+tmp[4224]*kernel[5]+tmp[4322]*kernel[6]+tmp[4323]*kernel[7]+tmp[4324]*kernel[8];
				ans[4224]<=tmp[4123]*kernel[0]+tmp[4124]*kernel[1]+tmp[4125]*kernel[2]+tmp[4223]*kernel[3]+tmp[4224]*kernel[4]+tmp[4225]*kernel[5]+tmp[4323]*kernel[6]+tmp[4324]*kernel[7]+tmp[4325]*kernel[8];
				ans[4225]<=tmp[4124]*kernel[0]+tmp[4125]*kernel[1]+tmp[4126]*kernel[2]+tmp[4224]*kernel[3]+tmp[4225]*kernel[4]+tmp[4226]*kernel[5]+tmp[4324]*kernel[6]+tmp[4325]*kernel[7]+tmp[4326]*kernel[8];
				ans[4226]<=tmp[4125]*kernel[0]+tmp[4126]*kernel[1]+tmp[4127]*kernel[2]+tmp[4225]*kernel[3]+tmp[4226]*kernel[4]+tmp[4227]*kernel[5]+tmp[4325]*kernel[6]+tmp[4326]*kernel[7]+tmp[4327]*kernel[8];
				ans[4227]<=tmp[4126]*kernel[0]+tmp[4127]*kernel[1]+tmp[4128]*kernel[2]+tmp[4226]*kernel[3]+tmp[4227]*kernel[4]+tmp[4228]*kernel[5]+tmp[4326]*kernel[6]+tmp[4327]*kernel[7]+tmp[4328]*kernel[8];
				ans[4228]<=tmp[4127]*kernel[0]+tmp[4128]*kernel[1]+tmp[4129]*kernel[2]+tmp[4227]*kernel[3]+tmp[4228]*kernel[4]+tmp[4229]*kernel[5]+tmp[4327]*kernel[6]+tmp[4328]*kernel[7]+tmp[4329]*kernel[8];
				ans[4229]<=tmp[4128]*kernel[0]+tmp[4129]*kernel[1]+tmp[4130]*kernel[2]+tmp[4228]*kernel[3]+tmp[4229]*kernel[4]+tmp[4230]*kernel[5]+tmp[4328]*kernel[6]+tmp[4329]*kernel[7]+tmp[4330]*kernel[8];
				ans[4230]<=tmp[4129]*kernel[0]+tmp[4130]*kernel[1]+tmp[4131]*kernel[2]+tmp[4229]*kernel[3]+tmp[4230]*kernel[4]+tmp[4231]*kernel[5]+tmp[4329]*kernel[6]+tmp[4330]*kernel[7]+tmp[4331]*kernel[8];
				ans[4231]<=tmp[4130]*kernel[0]+tmp[4131]*kernel[1]+tmp[4132]*kernel[2]+tmp[4230]*kernel[3]+tmp[4231]*kernel[4]+tmp[4232]*kernel[5]+tmp[4330]*kernel[6]+tmp[4331]*kernel[7]+tmp[4332]*kernel[8];
				ans[4232]<=tmp[4131]*kernel[0]+tmp[4132]*kernel[1]+tmp[4133]*kernel[2]+tmp[4231]*kernel[3]+tmp[4232]*kernel[4]+tmp[4233]*kernel[5]+tmp[4331]*kernel[6]+tmp[4332]*kernel[7]+tmp[4333]*kernel[8];
				ans[4233]<=tmp[4132]*kernel[0]+tmp[4133]*kernel[1]+tmp[4134]*kernel[2]+tmp[4232]*kernel[3]+tmp[4233]*kernel[4]+tmp[4234]*kernel[5]+tmp[4332]*kernel[6]+tmp[4333]*kernel[7]+tmp[4334]*kernel[8];
				ans[4234]<=tmp[4133]*kernel[0]+tmp[4134]*kernel[1]+tmp[4135]*kernel[2]+tmp[4233]*kernel[3]+tmp[4234]*kernel[4]+tmp[4235]*kernel[5]+tmp[4333]*kernel[6]+tmp[4334]*kernel[7]+tmp[4335]*kernel[8];
				ans[4235]<=tmp[4134]*kernel[0]+tmp[4135]*kernel[1]+tmp[4136]*kernel[2]+tmp[4234]*kernel[3]+tmp[4235]*kernel[4]+tmp[4236]*kernel[5]+tmp[4334]*kernel[6]+tmp[4335]*kernel[7]+tmp[4336]*kernel[8];
				ans[4236]<=tmp[4135]*kernel[0]+tmp[4136]*kernel[1]+tmp[4137]*kernel[2]+tmp[4235]*kernel[3]+tmp[4236]*kernel[4]+tmp[4237]*kernel[5]+tmp[4335]*kernel[6]+tmp[4336]*kernel[7]+tmp[4337]*kernel[8];
				ans[4237]<=tmp[4136]*kernel[0]+tmp[4137]*kernel[1]+tmp[4138]*kernel[2]+tmp[4236]*kernel[3]+tmp[4237]*kernel[4]+tmp[4238]*kernel[5]+tmp[4336]*kernel[6]+tmp[4337]*kernel[7]+tmp[4338]*kernel[8];
				ans[4238]<=tmp[4137]*kernel[0]+tmp[4138]*kernel[1]+tmp[4139]*kernel[2]+tmp[4237]*kernel[3]+tmp[4238]*kernel[4]+tmp[4239]*kernel[5]+tmp[4337]*kernel[6]+tmp[4338]*kernel[7]+tmp[4339]*kernel[8];
				ans[4239]<=tmp[4138]*kernel[0]+tmp[4139]*kernel[1]+tmp[4140]*kernel[2]+tmp[4238]*kernel[3]+tmp[4239]*kernel[4]+tmp[4240]*kernel[5]+tmp[4338]*kernel[6]+tmp[4339]*kernel[7]+tmp[4340]*kernel[8];
				ans[4240]<=tmp[4139]*kernel[0]+tmp[4140]*kernel[1]+tmp[4141]*kernel[2]+tmp[4239]*kernel[3]+tmp[4240]*kernel[4]+tmp[4241]*kernel[5]+tmp[4339]*kernel[6]+tmp[4340]*kernel[7]+tmp[4341]*kernel[8];
				ans[4241]<=tmp[4140]*kernel[0]+tmp[4141]*kernel[1]+tmp[4142]*kernel[2]+tmp[4240]*kernel[3]+tmp[4241]*kernel[4]+tmp[4242]*kernel[5]+tmp[4340]*kernel[6]+tmp[4341]*kernel[7]+tmp[4342]*kernel[8];
				ans[4242]<=tmp[4141]*kernel[0]+tmp[4142]*kernel[1]+tmp[4143]*kernel[2]+tmp[4241]*kernel[3]+tmp[4242]*kernel[4]+tmp[4243]*kernel[5]+tmp[4341]*kernel[6]+tmp[4342]*kernel[7]+tmp[4343]*kernel[8];
				ans[4243]<=tmp[4142]*kernel[0]+tmp[4143]*kernel[1]+tmp[4144]*kernel[2]+tmp[4242]*kernel[3]+tmp[4243]*kernel[4]+tmp[4244]*kernel[5]+tmp[4342]*kernel[6]+tmp[4343]*kernel[7]+tmp[4344]*kernel[8];
				ans[4244]<=tmp[4143]*kernel[0]+tmp[4144]*kernel[1]+tmp[4145]*kernel[2]+tmp[4243]*kernel[3]+tmp[4244]*kernel[4]+tmp[4245]*kernel[5]+tmp[4343]*kernel[6]+tmp[4344]*kernel[7]+tmp[4345]*kernel[8];
				ans[4245]<=tmp[4144]*kernel[0]+tmp[4145]*kernel[1]+tmp[4146]*kernel[2]+tmp[4244]*kernel[3]+tmp[4245]*kernel[4]+tmp[4246]*kernel[5]+tmp[4344]*kernel[6]+tmp[4345]*kernel[7]+tmp[4346]*kernel[8];
				ans[4246]<=tmp[4145]*kernel[0]+tmp[4146]*kernel[1]+tmp[4147]*kernel[2]+tmp[4245]*kernel[3]+tmp[4246]*kernel[4]+tmp[4247]*kernel[5]+tmp[4345]*kernel[6]+tmp[4346]*kernel[7]+tmp[4347]*kernel[8];
				ans[4247]<=tmp[4146]*kernel[0]+tmp[4147]*kernel[1]+tmp[4148]*kernel[2]+tmp[4246]*kernel[3]+tmp[4247]*kernel[4]+tmp[4248]*kernel[5]+tmp[4346]*kernel[6]+tmp[4347]*kernel[7]+tmp[4348]*kernel[8];
				ans[4248]<=tmp[4147]*kernel[0]+tmp[4148]*kernel[1]+tmp[4149]*kernel[2]+tmp[4247]*kernel[3]+tmp[4248]*kernel[4]+tmp[4249]*kernel[5]+tmp[4347]*kernel[6]+tmp[4348]*kernel[7]+tmp[4349]*kernel[8];
				ans[4249]<=tmp[4148]*kernel[0]+tmp[4149]*kernel[1]+tmp[4150]*kernel[2]+tmp[4248]*kernel[3]+tmp[4249]*kernel[4]+tmp[4250]*kernel[5]+tmp[4348]*kernel[6]+tmp[4349]*kernel[7]+tmp[4350]*kernel[8];
				ans[4250]<=tmp[4149]*kernel[0]+tmp[4150]*kernel[1]+tmp[4151]*kernel[2]+tmp[4249]*kernel[3]+tmp[4250]*kernel[4]+tmp[4251]*kernel[5]+tmp[4349]*kernel[6]+tmp[4350]*kernel[7]+tmp[4351]*kernel[8];
				ans[4251]<=tmp[4150]*kernel[0]+tmp[4151]*kernel[1]+tmp[4152]*kernel[2]+tmp[4250]*kernel[3]+tmp[4251]*kernel[4]+tmp[4252]*kernel[5]+tmp[4350]*kernel[6]+tmp[4351]*kernel[7]+tmp[4352]*kernel[8];
				ans[4252]<=tmp[4151]*kernel[0]+tmp[4152]*kernel[1]+tmp[4153]*kernel[2]+tmp[4251]*kernel[3]+tmp[4252]*kernel[4]+tmp[4253]*kernel[5]+tmp[4351]*kernel[6]+tmp[4352]*kernel[7]+tmp[4353]*kernel[8];
				ans[4253]<=tmp[4152]*kernel[0]+tmp[4153]*kernel[1]+tmp[4154]*kernel[2]+tmp[4252]*kernel[3]+tmp[4253]*kernel[4]+tmp[4254]*kernel[5]+tmp[4352]*kernel[6]+tmp[4353]*kernel[7]+tmp[4354]*kernel[8];
				ans[4254]<=tmp[4153]*kernel[0]+tmp[4154]*kernel[1]+tmp[4155]*kernel[2]+tmp[4253]*kernel[3]+tmp[4254]*kernel[4]+tmp[4255]*kernel[5]+tmp[4353]*kernel[6]+tmp[4354]*kernel[7]+tmp[4355]*kernel[8];
				ans[4255]<=tmp[4154]*kernel[0]+tmp[4155]*kernel[1]+tmp[4156]*kernel[2]+tmp[4254]*kernel[3]+tmp[4255]*kernel[4]+tmp[4256]*kernel[5]+tmp[4354]*kernel[6]+tmp[4355]*kernel[7]+tmp[4356]*kernel[8];
				ans[4256]<=tmp[4155]*kernel[0]+tmp[4156]*kernel[1]+tmp[4157]*kernel[2]+tmp[4255]*kernel[3]+tmp[4256]*kernel[4]+tmp[4257]*kernel[5]+tmp[4355]*kernel[6]+tmp[4356]*kernel[7]+tmp[4357]*kernel[8];
				ans[4257]<=tmp[4156]*kernel[0]+tmp[4157]*kernel[1]+tmp[4158]*kernel[2]+tmp[4256]*kernel[3]+tmp[4257]*kernel[4]+tmp[4258]*kernel[5]+tmp[4356]*kernel[6]+tmp[4357]*kernel[7]+tmp[4358]*kernel[8];
				ans[4258]<=tmp[4157]*kernel[0]+tmp[4158]*kernel[1]+tmp[4159]*kernel[2]+tmp[4257]*kernel[3]+tmp[4258]*kernel[4]+tmp[4259]*kernel[5]+tmp[4357]*kernel[6]+tmp[4358]*kernel[7]+tmp[4359]*kernel[8];
				ans[4259]<=tmp[4158]*kernel[0]+tmp[4159]*kernel[1]+tmp[4160]*kernel[2]+tmp[4258]*kernel[3]+tmp[4259]*kernel[4]+tmp[4260]*kernel[5]+tmp[4358]*kernel[6]+tmp[4359]*kernel[7]+tmp[4360]*kernel[8];
				ans[4260]<=tmp[4159]*kernel[0]+tmp[4160]*kernel[1]+tmp[4161]*kernel[2]+tmp[4259]*kernel[3]+tmp[4260]*kernel[4]+tmp[4261]*kernel[5]+tmp[4359]*kernel[6]+tmp[4360]*kernel[7]+tmp[4361]*kernel[8];
				ans[4261]<=tmp[4160]*kernel[0]+tmp[4161]*kernel[1]+tmp[4162]*kernel[2]+tmp[4260]*kernel[3]+tmp[4261]*kernel[4]+tmp[4262]*kernel[5]+tmp[4360]*kernel[6]+tmp[4361]*kernel[7]+tmp[4362]*kernel[8];
				ans[4262]<=tmp[4161]*kernel[0]+tmp[4162]*kernel[1]+tmp[4163]*kernel[2]+tmp[4261]*kernel[3]+tmp[4262]*kernel[4]+tmp[4263]*kernel[5]+tmp[4361]*kernel[6]+tmp[4362]*kernel[7]+tmp[4363]*kernel[8];
				ans[4263]<=tmp[4162]*kernel[0]+tmp[4163]*kernel[1]+tmp[4164]*kernel[2]+tmp[4262]*kernel[3]+tmp[4263]*kernel[4]+tmp[4264]*kernel[5]+tmp[4362]*kernel[6]+tmp[4363]*kernel[7]+tmp[4364]*kernel[8];
				ans[4264]<=tmp[4163]*kernel[0]+tmp[4164]*kernel[1]+tmp[4165]*kernel[2]+tmp[4263]*kernel[3]+tmp[4264]*kernel[4]+tmp[4265]*kernel[5]+tmp[4363]*kernel[6]+tmp[4364]*kernel[7]+tmp[4365]*kernel[8];
				ans[4265]<=tmp[4164]*kernel[0]+tmp[4165]*kernel[1]+tmp[4166]*kernel[2]+tmp[4264]*kernel[3]+tmp[4265]*kernel[4]+tmp[4266]*kernel[5]+tmp[4364]*kernel[6]+tmp[4365]*kernel[7]+tmp[4366]*kernel[8];
				ans[4266]<=tmp[4165]*kernel[0]+tmp[4166]*kernel[1]+tmp[4167]*kernel[2]+tmp[4265]*kernel[3]+tmp[4266]*kernel[4]+tmp[4267]*kernel[5]+tmp[4365]*kernel[6]+tmp[4366]*kernel[7]+tmp[4367]*kernel[8];
				ans[4267]<=tmp[4166]*kernel[0]+tmp[4167]*kernel[1]+tmp[4168]*kernel[2]+tmp[4266]*kernel[3]+tmp[4267]*kernel[4]+tmp[4268]*kernel[5]+tmp[4366]*kernel[6]+tmp[4367]*kernel[7]+tmp[4368]*kernel[8];
				ans[4268]<=tmp[4167]*kernel[0]+tmp[4168]*kernel[1]+tmp[4169]*kernel[2]+tmp[4267]*kernel[3]+tmp[4268]*kernel[4]+tmp[4269]*kernel[5]+tmp[4367]*kernel[6]+tmp[4368]*kernel[7]+tmp[4369]*kernel[8];
				ans[4269]<=tmp[4168]*kernel[0]+tmp[4169]*kernel[1]+tmp[4170]*kernel[2]+tmp[4268]*kernel[3]+tmp[4269]*kernel[4]+tmp[4270]*kernel[5]+tmp[4368]*kernel[6]+tmp[4369]*kernel[7]+tmp[4370]*kernel[8];
				ans[4270]<=tmp[4169]*kernel[0]+tmp[4170]*kernel[1]+tmp[4171]*kernel[2]+tmp[4269]*kernel[3]+tmp[4270]*kernel[4]+tmp[4271]*kernel[5]+tmp[4369]*kernel[6]+tmp[4370]*kernel[7]+tmp[4371]*kernel[8];
				ans[4271]<=tmp[4170]*kernel[0]+tmp[4171]*kernel[1]+tmp[4172]*kernel[2]+tmp[4270]*kernel[3]+tmp[4271]*kernel[4]+tmp[4272]*kernel[5]+tmp[4370]*kernel[6]+tmp[4371]*kernel[7]+tmp[4372]*kernel[8];
				ans[4272]<=tmp[4171]*kernel[0]+tmp[4172]*kernel[1]+tmp[4173]*kernel[2]+tmp[4271]*kernel[3]+tmp[4272]*kernel[4]+tmp[4273]*kernel[5]+tmp[4371]*kernel[6]+tmp[4372]*kernel[7]+tmp[4373]*kernel[8];
				ans[4273]<=tmp[4172]*kernel[0]+tmp[4173]*kernel[1]+tmp[4174]*kernel[2]+tmp[4272]*kernel[3]+tmp[4273]*kernel[4]+tmp[4274]*kernel[5]+tmp[4372]*kernel[6]+tmp[4373]*kernel[7]+tmp[4374]*kernel[8];
				ans[4274]<=tmp[4173]*kernel[0]+tmp[4174]*kernel[1]+tmp[4175]*kernel[2]+tmp[4273]*kernel[3]+tmp[4274]*kernel[4]+tmp[4275]*kernel[5]+tmp[4373]*kernel[6]+tmp[4374]*kernel[7]+tmp[4375]*kernel[8];
				ans[4275]<=tmp[4174]*kernel[0]+tmp[4175]*kernel[1]+tmp[4176]*kernel[2]+tmp[4274]*kernel[3]+tmp[4275]*kernel[4]+tmp[4276]*kernel[5]+tmp[4374]*kernel[6]+tmp[4375]*kernel[7]+tmp[4376]*kernel[8];
				ans[4276]<=tmp[4175]*kernel[0]+tmp[4176]*kernel[1]+tmp[4177]*kernel[2]+tmp[4275]*kernel[3]+tmp[4276]*kernel[4]+tmp[4277]*kernel[5]+tmp[4375]*kernel[6]+tmp[4376]*kernel[7]+tmp[4377]*kernel[8];
				ans[4277]<=tmp[4176]*kernel[0]+tmp[4177]*kernel[1]+tmp[4178]*kernel[2]+tmp[4276]*kernel[3]+tmp[4277]*kernel[4]+tmp[4278]*kernel[5]+tmp[4376]*kernel[6]+tmp[4377]*kernel[7]+tmp[4378]*kernel[8];
				ans[4278]<=tmp[4177]*kernel[0]+tmp[4178]*kernel[1]+tmp[4179]*kernel[2]+tmp[4277]*kernel[3]+tmp[4278]*kernel[4]+tmp[4279]*kernel[5]+tmp[4377]*kernel[6]+tmp[4378]*kernel[7]+tmp[4379]*kernel[8];
				ans[4279]<=tmp[4178]*kernel[0]+tmp[4179]*kernel[1]+tmp[4180]*kernel[2]+tmp[4278]*kernel[3]+tmp[4279]*kernel[4]+tmp[4280]*kernel[5]+tmp[4378]*kernel[6]+tmp[4379]*kernel[7]+tmp[4380]*kernel[8];
				ans[4280]<=tmp[4179]*kernel[0]+tmp[4180]*kernel[1]+tmp[4181]*kernel[2]+tmp[4279]*kernel[3]+tmp[4280]*kernel[4]+tmp[4281]*kernel[5]+tmp[4379]*kernel[6]+tmp[4380]*kernel[7]+tmp[4381]*kernel[8];
				ans[4281]<=tmp[4180]*kernel[0]+tmp[4181]*kernel[1]+tmp[4182]*kernel[2]+tmp[4280]*kernel[3]+tmp[4281]*kernel[4]+tmp[4282]*kernel[5]+tmp[4380]*kernel[6]+tmp[4381]*kernel[7]+tmp[4382]*kernel[8];
				ans[4282]<=tmp[4181]*kernel[0]+tmp[4182]*kernel[1]+tmp[4183]*kernel[2]+tmp[4281]*kernel[3]+tmp[4282]*kernel[4]+tmp[4283]*kernel[5]+tmp[4381]*kernel[6]+tmp[4382]*kernel[7]+tmp[4383]*kernel[8];
				ans[4283]<=tmp[4182]*kernel[0]+tmp[4183]*kernel[1]+tmp[4184]*kernel[2]+tmp[4282]*kernel[3]+tmp[4283]*kernel[4]+tmp[4284]*kernel[5]+tmp[4382]*kernel[6]+tmp[4383]*kernel[7]+tmp[4384]*kernel[8];
				ans[4284]<=tmp[4183]*kernel[0]+tmp[4184]*kernel[1]+tmp[4185]*kernel[2]+tmp[4283]*kernel[3]+tmp[4284]*kernel[4]+tmp[4285]*kernel[5]+tmp[4383]*kernel[6]+tmp[4384]*kernel[7]+tmp[4385]*kernel[8];
				ans[4285]<=tmp[4184]*kernel[0]+tmp[4185]*kernel[1]+tmp[4186]*kernel[2]+tmp[4284]*kernel[3]+tmp[4285]*kernel[4]+tmp[4286]*kernel[5]+tmp[4384]*kernel[6]+tmp[4385]*kernel[7]+tmp[4386]*kernel[8];
				ans[4286]<=tmp[4185]*kernel[0]+tmp[4186]*kernel[1]+tmp[4187]*kernel[2]+tmp[4285]*kernel[3]+tmp[4286]*kernel[4]+tmp[4287]*kernel[5]+tmp[4385]*kernel[6]+tmp[4386]*kernel[7]+tmp[4387]*kernel[8];
				ans[4287]<=tmp[4186]*kernel[0]+tmp[4187]*kernel[1]+tmp[4188]*kernel[2]+tmp[4286]*kernel[3]+tmp[4287]*kernel[4]+tmp[4288]*kernel[5]+tmp[4386]*kernel[6]+tmp[4387]*kernel[7]+tmp[4388]*kernel[8];
				ans[4288]<=tmp[4187]*kernel[0]+tmp[4188]*kernel[1]+tmp[4189]*kernel[2]+tmp[4287]*kernel[3]+tmp[4288]*kernel[4]+tmp[4289]*kernel[5]+tmp[4387]*kernel[6]+tmp[4388]*kernel[7]+tmp[4389]*kernel[8];
				ans[4289]<=tmp[4188]*kernel[0]+tmp[4189]*kernel[1]+tmp[4190]*kernel[2]+tmp[4288]*kernel[3]+tmp[4289]*kernel[4]+tmp[4290]*kernel[5]+tmp[4388]*kernel[6]+tmp[4389]*kernel[7]+tmp[4390]*kernel[8];
				ans[4290]<=tmp[4189]*kernel[0]+tmp[4190]*kernel[1]+tmp[4191]*kernel[2]+tmp[4289]*kernel[3]+tmp[4290]*kernel[4]+tmp[4291]*kernel[5]+tmp[4389]*kernel[6]+tmp[4390]*kernel[7]+tmp[4391]*kernel[8];
				ans[4291]<=tmp[4190]*kernel[0]+tmp[4191]*kernel[1]+tmp[4192]*kernel[2]+tmp[4290]*kernel[3]+tmp[4291]*kernel[4]+tmp[4292]*kernel[5]+tmp[4390]*kernel[6]+tmp[4391]*kernel[7]+tmp[4392]*kernel[8];
				ans[4292]<=tmp[4191]*kernel[0]+tmp[4192]*kernel[1]+tmp[4193]*kernel[2]+tmp[4291]*kernel[3]+tmp[4292]*kernel[4]+tmp[4293]*kernel[5]+tmp[4391]*kernel[6]+tmp[4392]*kernel[7]+tmp[4393]*kernel[8];
				ans[4293]<=tmp[4192]*kernel[0]+tmp[4193]*kernel[1]+tmp[4194]*kernel[2]+tmp[4292]*kernel[3]+tmp[4293]*kernel[4]+tmp[4294]*kernel[5]+tmp[4392]*kernel[6]+tmp[4393]*kernel[7]+tmp[4394]*kernel[8];
				ans[4294]<=tmp[4193]*kernel[0]+tmp[4194]*kernel[1]+tmp[4195]*kernel[2]+tmp[4293]*kernel[3]+tmp[4294]*kernel[4]+tmp[4295]*kernel[5]+tmp[4393]*kernel[6]+tmp[4394]*kernel[7]+tmp[4395]*kernel[8];
				ans[4295]<=tmp[4194]*kernel[0]+tmp[4195]*kernel[1]+tmp[4196]*kernel[2]+tmp[4294]*kernel[3]+tmp[4295]*kernel[4]+tmp[4296]*kernel[5]+tmp[4394]*kernel[6]+tmp[4395]*kernel[7]+tmp[4396]*kernel[8];
				ans[4296]<=tmp[4195]*kernel[0]+tmp[4196]*kernel[1]+tmp[4197]*kernel[2]+tmp[4295]*kernel[3]+tmp[4296]*kernel[4]+tmp[4297]*kernel[5]+tmp[4395]*kernel[6]+tmp[4396]*kernel[7]+tmp[4397]*kernel[8];
				ans[4297]<=tmp[4196]*kernel[0]+tmp[4197]*kernel[1]+tmp[4198]*kernel[2]+tmp[4296]*kernel[3]+tmp[4297]*kernel[4]+tmp[4298]*kernel[5]+tmp[4396]*kernel[6]+tmp[4397]*kernel[7]+tmp[4398]*kernel[8];
				ans[4298]<=tmp[4197]*kernel[0]+tmp[4198]*kernel[1]+tmp[4199]*kernel[2]+tmp[4297]*kernel[3]+tmp[4298]*kernel[4]+tmp[4299]*kernel[5]+tmp[4397]*kernel[6]+tmp[4398]*kernel[7]+tmp[4399]*kernel[8];
				ans[4299]<=tmp[4198]*kernel[0]+tmp[4199]*kernel[1]+tmp[4298]*kernel[3]+tmp[4299]*kernel[4]+tmp[4398]*kernel[6]+tmp[4399]*kernel[7];
				ans[4300]<=tmp[4200]*kernel[1]+tmp[4201]*kernel[2]+tmp[4300]*kernel[4]+tmp[4301]*kernel[5]+tmp[4400]*kernel[7]+tmp[4401]*kernel[8];
				ans[4301]<=tmp[4200]*kernel[0]+tmp[4201]*kernel[1]+tmp[4202]*kernel[2]+tmp[4300]*kernel[3]+tmp[4301]*kernel[4]+tmp[4302]*kernel[5]+tmp[4400]*kernel[6]+tmp[4401]*kernel[7]+tmp[4402]*kernel[8];
				ans[4302]<=tmp[4201]*kernel[0]+tmp[4202]*kernel[1]+tmp[4203]*kernel[2]+tmp[4301]*kernel[3]+tmp[4302]*kernel[4]+tmp[4303]*kernel[5]+tmp[4401]*kernel[6]+tmp[4402]*kernel[7]+tmp[4403]*kernel[8];
				ans[4303]<=tmp[4202]*kernel[0]+tmp[4203]*kernel[1]+tmp[4204]*kernel[2]+tmp[4302]*kernel[3]+tmp[4303]*kernel[4]+tmp[4304]*kernel[5]+tmp[4402]*kernel[6]+tmp[4403]*kernel[7]+tmp[4404]*kernel[8];
				ans[4304]<=tmp[4203]*kernel[0]+tmp[4204]*kernel[1]+tmp[4205]*kernel[2]+tmp[4303]*kernel[3]+tmp[4304]*kernel[4]+tmp[4305]*kernel[5]+tmp[4403]*kernel[6]+tmp[4404]*kernel[7]+tmp[4405]*kernel[8];
				ans[4305]<=tmp[4204]*kernel[0]+tmp[4205]*kernel[1]+tmp[4206]*kernel[2]+tmp[4304]*kernel[3]+tmp[4305]*kernel[4]+tmp[4306]*kernel[5]+tmp[4404]*kernel[6]+tmp[4405]*kernel[7]+tmp[4406]*kernel[8];
				ans[4306]<=tmp[4205]*kernel[0]+tmp[4206]*kernel[1]+tmp[4207]*kernel[2]+tmp[4305]*kernel[3]+tmp[4306]*kernel[4]+tmp[4307]*kernel[5]+tmp[4405]*kernel[6]+tmp[4406]*kernel[7]+tmp[4407]*kernel[8];
				ans[4307]<=tmp[4206]*kernel[0]+tmp[4207]*kernel[1]+tmp[4208]*kernel[2]+tmp[4306]*kernel[3]+tmp[4307]*kernel[4]+tmp[4308]*kernel[5]+tmp[4406]*kernel[6]+tmp[4407]*kernel[7]+tmp[4408]*kernel[8];
				ans[4308]<=tmp[4207]*kernel[0]+tmp[4208]*kernel[1]+tmp[4209]*kernel[2]+tmp[4307]*kernel[3]+tmp[4308]*kernel[4]+tmp[4309]*kernel[5]+tmp[4407]*kernel[6]+tmp[4408]*kernel[7]+tmp[4409]*kernel[8];
				ans[4309]<=tmp[4208]*kernel[0]+tmp[4209]*kernel[1]+tmp[4210]*kernel[2]+tmp[4308]*kernel[3]+tmp[4309]*kernel[4]+tmp[4310]*kernel[5]+tmp[4408]*kernel[6]+tmp[4409]*kernel[7]+tmp[4410]*kernel[8];
				ans[4310]<=tmp[4209]*kernel[0]+tmp[4210]*kernel[1]+tmp[4211]*kernel[2]+tmp[4309]*kernel[3]+tmp[4310]*kernel[4]+tmp[4311]*kernel[5]+tmp[4409]*kernel[6]+tmp[4410]*kernel[7]+tmp[4411]*kernel[8];
				ans[4311]<=tmp[4210]*kernel[0]+tmp[4211]*kernel[1]+tmp[4212]*kernel[2]+tmp[4310]*kernel[3]+tmp[4311]*kernel[4]+tmp[4312]*kernel[5]+tmp[4410]*kernel[6]+tmp[4411]*kernel[7]+tmp[4412]*kernel[8];
				ans[4312]<=tmp[4211]*kernel[0]+tmp[4212]*kernel[1]+tmp[4213]*kernel[2]+tmp[4311]*kernel[3]+tmp[4312]*kernel[4]+tmp[4313]*kernel[5]+tmp[4411]*kernel[6]+tmp[4412]*kernel[7]+tmp[4413]*kernel[8];
				ans[4313]<=tmp[4212]*kernel[0]+tmp[4213]*kernel[1]+tmp[4214]*kernel[2]+tmp[4312]*kernel[3]+tmp[4313]*kernel[4]+tmp[4314]*kernel[5]+tmp[4412]*kernel[6]+tmp[4413]*kernel[7]+tmp[4414]*kernel[8];
				ans[4314]<=tmp[4213]*kernel[0]+tmp[4214]*kernel[1]+tmp[4215]*kernel[2]+tmp[4313]*kernel[3]+tmp[4314]*kernel[4]+tmp[4315]*kernel[5]+tmp[4413]*kernel[6]+tmp[4414]*kernel[7]+tmp[4415]*kernel[8];
				ans[4315]<=tmp[4214]*kernel[0]+tmp[4215]*kernel[1]+tmp[4216]*kernel[2]+tmp[4314]*kernel[3]+tmp[4315]*kernel[4]+tmp[4316]*kernel[5]+tmp[4414]*kernel[6]+tmp[4415]*kernel[7]+tmp[4416]*kernel[8];
				ans[4316]<=tmp[4215]*kernel[0]+tmp[4216]*kernel[1]+tmp[4217]*kernel[2]+tmp[4315]*kernel[3]+tmp[4316]*kernel[4]+tmp[4317]*kernel[5]+tmp[4415]*kernel[6]+tmp[4416]*kernel[7]+tmp[4417]*kernel[8];
				ans[4317]<=tmp[4216]*kernel[0]+tmp[4217]*kernel[1]+tmp[4218]*kernel[2]+tmp[4316]*kernel[3]+tmp[4317]*kernel[4]+tmp[4318]*kernel[5]+tmp[4416]*kernel[6]+tmp[4417]*kernel[7]+tmp[4418]*kernel[8];
				ans[4318]<=tmp[4217]*kernel[0]+tmp[4218]*kernel[1]+tmp[4219]*kernel[2]+tmp[4317]*kernel[3]+tmp[4318]*kernel[4]+tmp[4319]*kernel[5]+tmp[4417]*kernel[6]+tmp[4418]*kernel[7]+tmp[4419]*kernel[8];
				ans[4319]<=tmp[4218]*kernel[0]+tmp[4219]*kernel[1]+tmp[4220]*kernel[2]+tmp[4318]*kernel[3]+tmp[4319]*kernel[4]+tmp[4320]*kernel[5]+tmp[4418]*kernel[6]+tmp[4419]*kernel[7]+tmp[4420]*kernel[8];
				ans[4320]<=tmp[4219]*kernel[0]+tmp[4220]*kernel[1]+tmp[4221]*kernel[2]+tmp[4319]*kernel[3]+tmp[4320]*kernel[4]+tmp[4321]*kernel[5]+tmp[4419]*kernel[6]+tmp[4420]*kernel[7]+tmp[4421]*kernel[8];
				ans[4321]<=tmp[4220]*kernel[0]+tmp[4221]*kernel[1]+tmp[4222]*kernel[2]+tmp[4320]*kernel[3]+tmp[4321]*kernel[4]+tmp[4322]*kernel[5]+tmp[4420]*kernel[6]+tmp[4421]*kernel[7]+tmp[4422]*kernel[8];
				ans[4322]<=tmp[4221]*kernel[0]+tmp[4222]*kernel[1]+tmp[4223]*kernel[2]+tmp[4321]*kernel[3]+tmp[4322]*kernel[4]+tmp[4323]*kernel[5]+tmp[4421]*kernel[6]+tmp[4422]*kernel[7]+tmp[4423]*kernel[8];
				ans[4323]<=tmp[4222]*kernel[0]+tmp[4223]*kernel[1]+tmp[4224]*kernel[2]+tmp[4322]*kernel[3]+tmp[4323]*kernel[4]+tmp[4324]*kernel[5]+tmp[4422]*kernel[6]+tmp[4423]*kernel[7]+tmp[4424]*kernel[8];
				ans[4324]<=tmp[4223]*kernel[0]+tmp[4224]*kernel[1]+tmp[4225]*kernel[2]+tmp[4323]*kernel[3]+tmp[4324]*kernel[4]+tmp[4325]*kernel[5]+tmp[4423]*kernel[6]+tmp[4424]*kernel[7]+tmp[4425]*kernel[8];
				ans[4325]<=tmp[4224]*kernel[0]+tmp[4225]*kernel[1]+tmp[4226]*kernel[2]+tmp[4324]*kernel[3]+tmp[4325]*kernel[4]+tmp[4326]*kernel[5]+tmp[4424]*kernel[6]+tmp[4425]*kernel[7]+tmp[4426]*kernel[8];
				ans[4326]<=tmp[4225]*kernel[0]+tmp[4226]*kernel[1]+tmp[4227]*kernel[2]+tmp[4325]*kernel[3]+tmp[4326]*kernel[4]+tmp[4327]*kernel[5]+tmp[4425]*kernel[6]+tmp[4426]*kernel[7]+tmp[4427]*kernel[8];
				ans[4327]<=tmp[4226]*kernel[0]+tmp[4227]*kernel[1]+tmp[4228]*kernel[2]+tmp[4326]*kernel[3]+tmp[4327]*kernel[4]+tmp[4328]*kernel[5]+tmp[4426]*kernel[6]+tmp[4427]*kernel[7]+tmp[4428]*kernel[8];
				ans[4328]<=tmp[4227]*kernel[0]+tmp[4228]*kernel[1]+tmp[4229]*kernel[2]+tmp[4327]*kernel[3]+tmp[4328]*kernel[4]+tmp[4329]*kernel[5]+tmp[4427]*kernel[6]+tmp[4428]*kernel[7]+tmp[4429]*kernel[8];
				ans[4329]<=tmp[4228]*kernel[0]+tmp[4229]*kernel[1]+tmp[4230]*kernel[2]+tmp[4328]*kernel[3]+tmp[4329]*kernel[4]+tmp[4330]*kernel[5]+tmp[4428]*kernel[6]+tmp[4429]*kernel[7]+tmp[4430]*kernel[8];
				ans[4330]<=tmp[4229]*kernel[0]+tmp[4230]*kernel[1]+tmp[4231]*kernel[2]+tmp[4329]*kernel[3]+tmp[4330]*kernel[4]+tmp[4331]*kernel[5]+tmp[4429]*kernel[6]+tmp[4430]*kernel[7]+tmp[4431]*kernel[8];
				ans[4331]<=tmp[4230]*kernel[0]+tmp[4231]*kernel[1]+tmp[4232]*kernel[2]+tmp[4330]*kernel[3]+tmp[4331]*kernel[4]+tmp[4332]*kernel[5]+tmp[4430]*kernel[6]+tmp[4431]*kernel[7]+tmp[4432]*kernel[8];
				ans[4332]<=tmp[4231]*kernel[0]+tmp[4232]*kernel[1]+tmp[4233]*kernel[2]+tmp[4331]*kernel[3]+tmp[4332]*kernel[4]+tmp[4333]*kernel[5]+tmp[4431]*kernel[6]+tmp[4432]*kernel[7]+tmp[4433]*kernel[8];
				ans[4333]<=tmp[4232]*kernel[0]+tmp[4233]*kernel[1]+tmp[4234]*kernel[2]+tmp[4332]*kernel[3]+tmp[4333]*kernel[4]+tmp[4334]*kernel[5]+tmp[4432]*kernel[6]+tmp[4433]*kernel[7]+tmp[4434]*kernel[8];
				ans[4334]<=tmp[4233]*kernel[0]+tmp[4234]*kernel[1]+tmp[4235]*kernel[2]+tmp[4333]*kernel[3]+tmp[4334]*kernel[4]+tmp[4335]*kernel[5]+tmp[4433]*kernel[6]+tmp[4434]*kernel[7]+tmp[4435]*kernel[8];
				ans[4335]<=tmp[4234]*kernel[0]+tmp[4235]*kernel[1]+tmp[4236]*kernel[2]+tmp[4334]*kernel[3]+tmp[4335]*kernel[4]+tmp[4336]*kernel[5]+tmp[4434]*kernel[6]+tmp[4435]*kernel[7]+tmp[4436]*kernel[8];
				ans[4336]<=tmp[4235]*kernel[0]+tmp[4236]*kernel[1]+tmp[4237]*kernel[2]+tmp[4335]*kernel[3]+tmp[4336]*kernel[4]+tmp[4337]*kernel[5]+tmp[4435]*kernel[6]+tmp[4436]*kernel[7]+tmp[4437]*kernel[8];
				ans[4337]<=tmp[4236]*kernel[0]+tmp[4237]*kernel[1]+tmp[4238]*kernel[2]+tmp[4336]*kernel[3]+tmp[4337]*kernel[4]+tmp[4338]*kernel[5]+tmp[4436]*kernel[6]+tmp[4437]*kernel[7]+tmp[4438]*kernel[8];
				ans[4338]<=tmp[4237]*kernel[0]+tmp[4238]*kernel[1]+tmp[4239]*kernel[2]+tmp[4337]*kernel[3]+tmp[4338]*kernel[4]+tmp[4339]*kernel[5]+tmp[4437]*kernel[6]+tmp[4438]*kernel[7]+tmp[4439]*kernel[8];
				ans[4339]<=tmp[4238]*kernel[0]+tmp[4239]*kernel[1]+tmp[4240]*kernel[2]+tmp[4338]*kernel[3]+tmp[4339]*kernel[4]+tmp[4340]*kernel[5]+tmp[4438]*kernel[6]+tmp[4439]*kernel[7]+tmp[4440]*kernel[8];
				ans[4340]<=tmp[4239]*kernel[0]+tmp[4240]*kernel[1]+tmp[4241]*kernel[2]+tmp[4339]*kernel[3]+tmp[4340]*kernel[4]+tmp[4341]*kernel[5]+tmp[4439]*kernel[6]+tmp[4440]*kernel[7]+tmp[4441]*kernel[8];
				ans[4341]<=tmp[4240]*kernel[0]+tmp[4241]*kernel[1]+tmp[4242]*kernel[2]+tmp[4340]*kernel[3]+tmp[4341]*kernel[4]+tmp[4342]*kernel[5]+tmp[4440]*kernel[6]+tmp[4441]*kernel[7]+tmp[4442]*kernel[8];
				ans[4342]<=tmp[4241]*kernel[0]+tmp[4242]*kernel[1]+tmp[4243]*kernel[2]+tmp[4341]*kernel[3]+tmp[4342]*kernel[4]+tmp[4343]*kernel[5]+tmp[4441]*kernel[6]+tmp[4442]*kernel[7]+tmp[4443]*kernel[8];
				ans[4343]<=tmp[4242]*kernel[0]+tmp[4243]*kernel[1]+tmp[4244]*kernel[2]+tmp[4342]*kernel[3]+tmp[4343]*kernel[4]+tmp[4344]*kernel[5]+tmp[4442]*kernel[6]+tmp[4443]*kernel[7]+tmp[4444]*kernel[8];
				ans[4344]<=tmp[4243]*kernel[0]+tmp[4244]*kernel[1]+tmp[4245]*kernel[2]+tmp[4343]*kernel[3]+tmp[4344]*kernel[4]+tmp[4345]*kernel[5]+tmp[4443]*kernel[6]+tmp[4444]*kernel[7]+tmp[4445]*kernel[8];
				ans[4345]<=tmp[4244]*kernel[0]+tmp[4245]*kernel[1]+tmp[4246]*kernel[2]+tmp[4344]*kernel[3]+tmp[4345]*kernel[4]+tmp[4346]*kernel[5]+tmp[4444]*kernel[6]+tmp[4445]*kernel[7]+tmp[4446]*kernel[8];
				ans[4346]<=tmp[4245]*kernel[0]+tmp[4246]*kernel[1]+tmp[4247]*kernel[2]+tmp[4345]*kernel[3]+tmp[4346]*kernel[4]+tmp[4347]*kernel[5]+tmp[4445]*kernel[6]+tmp[4446]*kernel[7]+tmp[4447]*kernel[8];
				ans[4347]<=tmp[4246]*kernel[0]+tmp[4247]*kernel[1]+tmp[4248]*kernel[2]+tmp[4346]*kernel[3]+tmp[4347]*kernel[4]+tmp[4348]*kernel[5]+tmp[4446]*kernel[6]+tmp[4447]*kernel[7]+tmp[4448]*kernel[8];
				ans[4348]<=tmp[4247]*kernel[0]+tmp[4248]*kernel[1]+tmp[4249]*kernel[2]+tmp[4347]*kernel[3]+tmp[4348]*kernel[4]+tmp[4349]*kernel[5]+tmp[4447]*kernel[6]+tmp[4448]*kernel[7]+tmp[4449]*kernel[8];
				ans[4349]<=tmp[4248]*kernel[0]+tmp[4249]*kernel[1]+tmp[4250]*kernel[2]+tmp[4348]*kernel[3]+tmp[4349]*kernel[4]+tmp[4350]*kernel[5]+tmp[4448]*kernel[6]+tmp[4449]*kernel[7]+tmp[4450]*kernel[8];
				ans[4350]<=tmp[4249]*kernel[0]+tmp[4250]*kernel[1]+tmp[4251]*kernel[2]+tmp[4349]*kernel[3]+tmp[4350]*kernel[4]+tmp[4351]*kernel[5]+tmp[4449]*kernel[6]+tmp[4450]*kernel[7]+tmp[4451]*kernel[8];
				ans[4351]<=tmp[4250]*kernel[0]+tmp[4251]*kernel[1]+tmp[4252]*kernel[2]+tmp[4350]*kernel[3]+tmp[4351]*kernel[4]+tmp[4352]*kernel[5]+tmp[4450]*kernel[6]+tmp[4451]*kernel[7]+tmp[4452]*kernel[8];
				ans[4352]<=tmp[4251]*kernel[0]+tmp[4252]*kernel[1]+tmp[4253]*kernel[2]+tmp[4351]*kernel[3]+tmp[4352]*kernel[4]+tmp[4353]*kernel[5]+tmp[4451]*kernel[6]+tmp[4452]*kernel[7]+tmp[4453]*kernel[8];
				ans[4353]<=tmp[4252]*kernel[0]+tmp[4253]*kernel[1]+tmp[4254]*kernel[2]+tmp[4352]*kernel[3]+tmp[4353]*kernel[4]+tmp[4354]*kernel[5]+tmp[4452]*kernel[6]+tmp[4453]*kernel[7]+tmp[4454]*kernel[8];
				ans[4354]<=tmp[4253]*kernel[0]+tmp[4254]*kernel[1]+tmp[4255]*kernel[2]+tmp[4353]*kernel[3]+tmp[4354]*kernel[4]+tmp[4355]*kernel[5]+tmp[4453]*kernel[6]+tmp[4454]*kernel[7]+tmp[4455]*kernel[8];
				ans[4355]<=tmp[4254]*kernel[0]+tmp[4255]*kernel[1]+tmp[4256]*kernel[2]+tmp[4354]*kernel[3]+tmp[4355]*kernel[4]+tmp[4356]*kernel[5]+tmp[4454]*kernel[6]+tmp[4455]*kernel[7]+tmp[4456]*kernel[8];
				ans[4356]<=tmp[4255]*kernel[0]+tmp[4256]*kernel[1]+tmp[4257]*kernel[2]+tmp[4355]*kernel[3]+tmp[4356]*kernel[4]+tmp[4357]*kernel[5]+tmp[4455]*kernel[6]+tmp[4456]*kernel[7]+tmp[4457]*kernel[8];
				ans[4357]<=tmp[4256]*kernel[0]+tmp[4257]*kernel[1]+tmp[4258]*kernel[2]+tmp[4356]*kernel[3]+tmp[4357]*kernel[4]+tmp[4358]*kernel[5]+tmp[4456]*kernel[6]+tmp[4457]*kernel[7]+tmp[4458]*kernel[8];
				ans[4358]<=tmp[4257]*kernel[0]+tmp[4258]*kernel[1]+tmp[4259]*kernel[2]+tmp[4357]*kernel[3]+tmp[4358]*kernel[4]+tmp[4359]*kernel[5]+tmp[4457]*kernel[6]+tmp[4458]*kernel[7]+tmp[4459]*kernel[8];
				ans[4359]<=tmp[4258]*kernel[0]+tmp[4259]*kernel[1]+tmp[4260]*kernel[2]+tmp[4358]*kernel[3]+tmp[4359]*kernel[4]+tmp[4360]*kernel[5]+tmp[4458]*kernel[6]+tmp[4459]*kernel[7]+tmp[4460]*kernel[8];
				ans[4360]<=tmp[4259]*kernel[0]+tmp[4260]*kernel[1]+tmp[4261]*kernel[2]+tmp[4359]*kernel[3]+tmp[4360]*kernel[4]+tmp[4361]*kernel[5]+tmp[4459]*kernel[6]+tmp[4460]*kernel[7]+tmp[4461]*kernel[8];
				ans[4361]<=tmp[4260]*kernel[0]+tmp[4261]*kernel[1]+tmp[4262]*kernel[2]+tmp[4360]*kernel[3]+tmp[4361]*kernel[4]+tmp[4362]*kernel[5]+tmp[4460]*kernel[6]+tmp[4461]*kernel[7]+tmp[4462]*kernel[8];
				ans[4362]<=tmp[4261]*kernel[0]+tmp[4262]*kernel[1]+tmp[4263]*kernel[2]+tmp[4361]*kernel[3]+tmp[4362]*kernel[4]+tmp[4363]*kernel[5]+tmp[4461]*kernel[6]+tmp[4462]*kernel[7]+tmp[4463]*kernel[8];
				ans[4363]<=tmp[4262]*kernel[0]+tmp[4263]*kernel[1]+tmp[4264]*kernel[2]+tmp[4362]*kernel[3]+tmp[4363]*kernel[4]+tmp[4364]*kernel[5]+tmp[4462]*kernel[6]+tmp[4463]*kernel[7]+tmp[4464]*kernel[8];
				ans[4364]<=tmp[4263]*kernel[0]+tmp[4264]*kernel[1]+tmp[4265]*kernel[2]+tmp[4363]*kernel[3]+tmp[4364]*kernel[4]+tmp[4365]*kernel[5]+tmp[4463]*kernel[6]+tmp[4464]*kernel[7]+tmp[4465]*kernel[8];
				ans[4365]<=tmp[4264]*kernel[0]+tmp[4265]*kernel[1]+tmp[4266]*kernel[2]+tmp[4364]*kernel[3]+tmp[4365]*kernel[4]+tmp[4366]*kernel[5]+tmp[4464]*kernel[6]+tmp[4465]*kernel[7]+tmp[4466]*kernel[8];
				ans[4366]<=tmp[4265]*kernel[0]+tmp[4266]*kernel[1]+tmp[4267]*kernel[2]+tmp[4365]*kernel[3]+tmp[4366]*kernel[4]+tmp[4367]*kernel[5]+tmp[4465]*kernel[6]+tmp[4466]*kernel[7]+tmp[4467]*kernel[8];
				ans[4367]<=tmp[4266]*kernel[0]+tmp[4267]*kernel[1]+tmp[4268]*kernel[2]+tmp[4366]*kernel[3]+tmp[4367]*kernel[4]+tmp[4368]*kernel[5]+tmp[4466]*kernel[6]+tmp[4467]*kernel[7]+tmp[4468]*kernel[8];
				ans[4368]<=tmp[4267]*kernel[0]+tmp[4268]*kernel[1]+tmp[4269]*kernel[2]+tmp[4367]*kernel[3]+tmp[4368]*kernel[4]+tmp[4369]*kernel[5]+tmp[4467]*kernel[6]+tmp[4468]*kernel[7]+tmp[4469]*kernel[8];
				ans[4369]<=tmp[4268]*kernel[0]+tmp[4269]*kernel[1]+tmp[4270]*kernel[2]+tmp[4368]*kernel[3]+tmp[4369]*kernel[4]+tmp[4370]*kernel[5]+tmp[4468]*kernel[6]+tmp[4469]*kernel[7]+tmp[4470]*kernel[8];
				ans[4370]<=tmp[4269]*kernel[0]+tmp[4270]*kernel[1]+tmp[4271]*kernel[2]+tmp[4369]*kernel[3]+tmp[4370]*kernel[4]+tmp[4371]*kernel[5]+tmp[4469]*kernel[6]+tmp[4470]*kernel[7]+tmp[4471]*kernel[8];
				ans[4371]<=tmp[4270]*kernel[0]+tmp[4271]*kernel[1]+tmp[4272]*kernel[2]+tmp[4370]*kernel[3]+tmp[4371]*kernel[4]+tmp[4372]*kernel[5]+tmp[4470]*kernel[6]+tmp[4471]*kernel[7]+tmp[4472]*kernel[8];
				ans[4372]<=tmp[4271]*kernel[0]+tmp[4272]*kernel[1]+tmp[4273]*kernel[2]+tmp[4371]*kernel[3]+tmp[4372]*kernel[4]+tmp[4373]*kernel[5]+tmp[4471]*kernel[6]+tmp[4472]*kernel[7]+tmp[4473]*kernel[8];
				ans[4373]<=tmp[4272]*kernel[0]+tmp[4273]*kernel[1]+tmp[4274]*kernel[2]+tmp[4372]*kernel[3]+tmp[4373]*kernel[4]+tmp[4374]*kernel[5]+tmp[4472]*kernel[6]+tmp[4473]*kernel[7]+tmp[4474]*kernel[8];
				ans[4374]<=tmp[4273]*kernel[0]+tmp[4274]*kernel[1]+tmp[4275]*kernel[2]+tmp[4373]*kernel[3]+tmp[4374]*kernel[4]+tmp[4375]*kernel[5]+tmp[4473]*kernel[6]+tmp[4474]*kernel[7]+tmp[4475]*kernel[8];
				ans[4375]<=tmp[4274]*kernel[0]+tmp[4275]*kernel[1]+tmp[4276]*kernel[2]+tmp[4374]*kernel[3]+tmp[4375]*kernel[4]+tmp[4376]*kernel[5]+tmp[4474]*kernel[6]+tmp[4475]*kernel[7]+tmp[4476]*kernel[8];
				ans[4376]<=tmp[4275]*kernel[0]+tmp[4276]*kernel[1]+tmp[4277]*kernel[2]+tmp[4375]*kernel[3]+tmp[4376]*kernel[4]+tmp[4377]*kernel[5]+tmp[4475]*kernel[6]+tmp[4476]*kernel[7]+tmp[4477]*kernel[8];
				ans[4377]<=tmp[4276]*kernel[0]+tmp[4277]*kernel[1]+tmp[4278]*kernel[2]+tmp[4376]*kernel[3]+tmp[4377]*kernel[4]+tmp[4378]*kernel[5]+tmp[4476]*kernel[6]+tmp[4477]*kernel[7]+tmp[4478]*kernel[8];
				ans[4378]<=tmp[4277]*kernel[0]+tmp[4278]*kernel[1]+tmp[4279]*kernel[2]+tmp[4377]*kernel[3]+tmp[4378]*kernel[4]+tmp[4379]*kernel[5]+tmp[4477]*kernel[6]+tmp[4478]*kernel[7]+tmp[4479]*kernel[8];
				ans[4379]<=tmp[4278]*kernel[0]+tmp[4279]*kernel[1]+tmp[4280]*kernel[2]+tmp[4378]*kernel[3]+tmp[4379]*kernel[4]+tmp[4380]*kernel[5]+tmp[4478]*kernel[6]+tmp[4479]*kernel[7]+tmp[4480]*kernel[8];
				ans[4380]<=tmp[4279]*kernel[0]+tmp[4280]*kernel[1]+tmp[4281]*kernel[2]+tmp[4379]*kernel[3]+tmp[4380]*kernel[4]+tmp[4381]*kernel[5]+tmp[4479]*kernel[6]+tmp[4480]*kernel[7]+tmp[4481]*kernel[8];
				ans[4381]<=tmp[4280]*kernel[0]+tmp[4281]*kernel[1]+tmp[4282]*kernel[2]+tmp[4380]*kernel[3]+tmp[4381]*kernel[4]+tmp[4382]*kernel[5]+tmp[4480]*kernel[6]+tmp[4481]*kernel[7]+tmp[4482]*kernel[8];
				ans[4382]<=tmp[4281]*kernel[0]+tmp[4282]*kernel[1]+tmp[4283]*kernel[2]+tmp[4381]*kernel[3]+tmp[4382]*kernel[4]+tmp[4383]*kernel[5]+tmp[4481]*kernel[6]+tmp[4482]*kernel[7]+tmp[4483]*kernel[8];
				ans[4383]<=tmp[4282]*kernel[0]+tmp[4283]*kernel[1]+tmp[4284]*kernel[2]+tmp[4382]*kernel[3]+tmp[4383]*kernel[4]+tmp[4384]*kernel[5]+tmp[4482]*kernel[6]+tmp[4483]*kernel[7]+tmp[4484]*kernel[8];
				ans[4384]<=tmp[4283]*kernel[0]+tmp[4284]*kernel[1]+tmp[4285]*kernel[2]+tmp[4383]*kernel[3]+tmp[4384]*kernel[4]+tmp[4385]*kernel[5]+tmp[4483]*kernel[6]+tmp[4484]*kernel[7]+tmp[4485]*kernel[8];
				ans[4385]<=tmp[4284]*kernel[0]+tmp[4285]*kernel[1]+tmp[4286]*kernel[2]+tmp[4384]*kernel[3]+tmp[4385]*kernel[4]+tmp[4386]*kernel[5]+tmp[4484]*kernel[6]+tmp[4485]*kernel[7]+tmp[4486]*kernel[8];
				ans[4386]<=tmp[4285]*kernel[0]+tmp[4286]*kernel[1]+tmp[4287]*kernel[2]+tmp[4385]*kernel[3]+tmp[4386]*kernel[4]+tmp[4387]*kernel[5]+tmp[4485]*kernel[6]+tmp[4486]*kernel[7]+tmp[4487]*kernel[8];
				ans[4387]<=tmp[4286]*kernel[0]+tmp[4287]*kernel[1]+tmp[4288]*kernel[2]+tmp[4386]*kernel[3]+tmp[4387]*kernel[4]+tmp[4388]*kernel[5]+tmp[4486]*kernel[6]+tmp[4487]*kernel[7]+tmp[4488]*kernel[8];
				ans[4388]<=tmp[4287]*kernel[0]+tmp[4288]*kernel[1]+tmp[4289]*kernel[2]+tmp[4387]*kernel[3]+tmp[4388]*kernel[4]+tmp[4389]*kernel[5]+tmp[4487]*kernel[6]+tmp[4488]*kernel[7]+tmp[4489]*kernel[8];
				ans[4389]<=tmp[4288]*kernel[0]+tmp[4289]*kernel[1]+tmp[4290]*kernel[2]+tmp[4388]*kernel[3]+tmp[4389]*kernel[4]+tmp[4390]*kernel[5]+tmp[4488]*kernel[6]+tmp[4489]*kernel[7]+tmp[4490]*kernel[8];
				ans[4390]<=tmp[4289]*kernel[0]+tmp[4290]*kernel[1]+tmp[4291]*kernel[2]+tmp[4389]*kernel[3]+tmp[4390]*kernel[4]+tmp[4391]*kernel[5]+tmp[4489]*kernel[6]+tmp[4490]*kernel[7]+tmp[4491]*kernel[8];
				ans[4391]<=tmp[4290]*kernel[0]+tmp[4291]*kernel[1]+tmp[4292]*kernel[2]+tmp[4390]*kernel[3]+tmp[4391]*kernel[4]+tmp[4392]*kernel[5]+tmp[4490]*kernel[6]+tmp[4491]*kernel[7]+tmp[4492]*kernel[8];
				ans[4392]<=tmp[4291]*kernel[0]+tmp[4292]*kernel[1]+tmp[4293]*kernel[2]+tmp[4391]*kernel[3]+tmp[4392]*kernel[4]+tmp[4393]*kernel[5]+tmp[4491]*kernel[6]+tmp[4492]*kernel[7]+tmp[4493]*kernel[8];
				ans[4393]<=tmp[4292]*kernel[0]+tmp[4293]*kernel[1]+tmp[4294]*kernel[2]+tmp[4392]*kernel[3]+tmp[4393]*kernel[4]+tmp[4394]*kernel[5]+tmp[4492]*kernel[6]+tmp[4493]*kernel[7]+tmp[4494]*kernel[8];
				ans[4394]<=tmp[4293]*kernel[0]+tmp[4294]*kernel[1]+tmp[4295]*kernel[2]+tmp[4393]*kernel[3]+tmp[4394]*kernel[4]+tmp[4395]*kernel[5]+tmp[4493]*kernel[6]+tmp[4494]*kernel[7]+tmp[4495]*kernel[8];
				ans[4395]<=tmp[4294]*kernel[0]+tmp[4295]*kernel[1]+tmp[4296]*kernel[2]+tmp[4394]*kernel[3]+tmp[4395]*kernel[4]+tmp[4396]*kernel[5]+tmp[4494]*kernel[6]+tmp[4495]*kernel[7]+tmp[4496]*kernel[8];
				ans[4396]<=tmp[4295]*kernel[0]+tmp[4296]*kernel[1]+tmp[4297]*kernel[2]+tmp[4395]*kernel[3]+tmp[4396]*kernel[4]+tmp[4397]*kernel[5]+tmp[4495]*kernel[6]+tmp[4496]*kernel[7]+tmp[4497]*kernel[8];
				ans[4397]<=tmp[4296]*kernel[0]+tmp[4297]*kernel[1]+tmp[4298]*kernel[2]+tmp[4396]*kernel[3]+tmp[4397]*kernel[4]+tmp[4398]*kernel[5]+tmp[4496]*kernel[6]+tmp[4497]*kernel[7]+tmp[4498]*kernel[8];
				ans[4398]<=tmp[4297]*kernel[0]+tmp[4298]*kernel[1]+tmp[4299]*kernel[2]+tmp[4397]*kernel[3]+tmp[4398]*kernel[4]+tmp[4399]*kernel[5]+tmp[4497]*kernel[6]+tmp[4498]*kernel[7]+tmp[4499]*kernel[8];
				ans[4399]<=tmp[4298]*kernel[0]+tmp[4299]*kernel[1]+tmp[4398]*kernel[3]+tmp[4399]*kernel[4]+tmp[4498]*kernel[6]+tmp[4499]*kernel[7];
				ans[4400]<=tmp[4300]*kernel[1]+tmp[4301]*kernel[2]+tmp[4400]*kernel[4]+tmp[4401]*kernel[5]+tmp[4500]*kernel[7]+tmp[4501]*kernel[8];
				ans[4401]<=tmp[4300]*kernel[0]+tmp[4301]*kernel[1]+tmp[4302]*kernel[2]+tmp[4400]*kernel[3]+tmp[4401]*kernel[4]+tmp[4402]*kernel[5]+tmp[4500]*kernel[6]+tmp[4501]*kernel[7]+tmp[4502]*kernel[8];
				ans[4402]<=tmp[4301]*kernel[0]+tmp[4302]*kernel[1]+tmp[4303]*kernel[2]+tmp[4401]*kernel[3]+tmp[4402]*kernel[4]+tmp[4403]*kernel[5]+tmp[4501]*kernel[6]+tmp[4502]*kernel[7]+tmp[4503]*kernel[8];
				ans[4403]<=tmp[4302]*kernel[0]+tmp[4303]*kernel[1]+tmp[4304]*kernel[2]+tmp[4402]*kernel[3]+tmp[4403]*kernel[4]+tmp[4404]*kernel[5]+tmp[4502]*kernel[6]+tmp[4503]*kernel[7]+tmp[4504]*kernel[8];
				ans[4404]<=tmp[4303]*kernel[0]+tmp[4304]*kernel[1]+tmp[4305]*kernel[2]+tmp[4403]*kernel[3]+tmp[4404]*kernel[4]+tmp[4405]*kernel[5]+tmp[4503]*kernel[6]+tmp[4504]*kernel[7]+tmp[4505]*kernel[8];
				ans[4405]<=tmp[4304]*kernel[0]+tmp[4305]*kernel[1]+tmp[4306]*kernel[2]+tmp[4404]*kernel[3]+tmp[4405]*kernel[4]+tmp[4406]*kernel[5]+tmp[4504]*kernel[6]+tmp[4505]*kernel[7]+tmp[4506]*kernel[8];
				ans[4406]<=tmp[4305]*kernel[0]+tmp[4306]*kernel[1]+tmp[4307]*kernel[2]+tmp[4405]*kernel[3]+tmp[4406]*kernel[4]+tmp[4407]*kernel[5]+tmp[4505]*kernel[6]+tmp[4506]*kernel[7]+tmp[4507]*kernel[8];
				ans[4407]<=tmp[4306]*kernel[0]+tmp[4307]*kernel[1]+tmp[4308]*kernel[2]+tmp[4406]*kernel[3]+tmp[4407]*kernel[4]+tmp[4408]*kernel[5]+tmp[4506]*kernel[6]+tmp[4507]*kernel[7]+tmp[4508]*kernel[8];
				ans[4408]<=tmp[4307]*kernel[0]+tmp[4308]*kernel[1]+tmp[4309]*kernel[2]+tmp[4407]*kernel[3]+tmp[4408]*kernel[4]+tmp[4409]*kernel[5]+tmp[4507]*kernel[6]+tmp[4508]*kernel[7]+tmp[4509]*kernel[8];
				ans[4409]<=tmp[4308]*kernel[0]+tmp[4309]*kernel[1]+tmp[4310]*kernel[2]+tmp[4408]*kernel[3]+tmp[4409]*kernel[4]+tmp[4410]*kernel[5]+tmp[4508]*kernel[6]+tmp[4509]*kernel[7]+tmp[4510]*kernel[8];
				ans[4410]<=tmp[4309]*kernel[0]+tmp[4310]*kernel[1]+tmp[4311]*kernel[2]+tmp[4409]*kernel[3]+tmp[4410]*kernel[4]+tmp[4411]*kernel[5]+tmp[4509]*kernel[6]+tmp[4510]*kernel[7]+tmp[4511]*kernel[8];
				ans[4411]<=tmp[4310]*kernel[0]+tmp[4311]*kernel[1]+tmp[4312]*kernel[2]+tmp[4410]*kernel[3]+tmp[4411]*kernel[4]+tmp[4412]*kernel[5]+tmp[4510]*kernel[6]+tmp[4511]*kernel[7]+tmp[4512]*kernel[8];
				ans[4412]<=tmp[4311]*kernel[0]+tmp[4312]*kernel[1]+tmp[4313]*kernel[2]+tmp[4411]*kernel[3]+tmp[4412]*kernel[4]+tmp[4413]*kernel[5]+tmp[4511]*kernel[6]+tmp[4512]*kernel[7]+tmp[4513]*kernel[8];
				ans[4413]<=tmp[4312]*kernel[0]+tmp[4313]*kernel[1]+tmp[4314]*kernel[2]+tmp[4412]*kernel[3]+tmp[4413]*kernel[4]+tmp[4414]*kernel[5]+tmp[4512]*kernel[6]+tmp[4513]*kernel[7]+tmp[4514]*kernel[8];
				ans[4414]<=tmp[4313]*kernel[0]+tmp[4314]*kernel[1]+tmp[4315]*kernel[2]+tmp[4413]*kernel[3]+tmp[4414]*kernel[4]+tmp[4415]*kernel[5]+tmp[4513]*kernel[6]+tmp[4514]*kernel[7]+tmp[4515]*kernel[8];
				ans[4415]<=tmp[4314]*kernel[0]+tmp[4315]*kernel[1]+tmp[4316]*kernel[2]+tmp[4414]*kernel[3]+tmp[4415]*kernel[4]+tmp[4416]*kernel[5]+tmp[4514]*kernel[6]+tmp[4515]*kernel[7]+tmp[4516]*kernel[8];
				ans[4416]<=tmp[4315]*kernel[0]+tmp[4316]*kernel[1]+tmp[4317]*kernel[2]+tmp[4415]*kernel[3]+tmp[4416]*kernel[4]+tmp[4417]*kernel[5]+tmp[4515]*kernel[6]+tmp[4516]*kernel[7]+tmp[4517]*kernel[8];
				ans[4417]<=tmp[4316]*kernel[0]+tmp[4317]*kernel[1]+tmp[4318]*kernel[2]+tmp[4416]*kernel[3]+tmp[4417]*kernel[4]+tmp[4418]*kernel[5]+tmp[4516]*kernel[6]+tmp[4517]*kernel[7]+tmp[4518]*kernel[8];
				ans[4418]<=tmp[4317]*kernel[0]+tmp[4318]*kernel[1]+tmp[4319]*kernel[2]+tmp[4417]*kernel[3]+tmp[4418]*kernel[4]+tmp[4419]*kernel[5]+tmp[4517]*kernel[6]+tmp[4518]*kernel[7]+tmp[4519]*kernel[8];
				ans[4419]<=tmp[4318]*kernel[0]+tmp[4319]*kernel[1]+tmp[4320]*kernel[2]+tmp[4418]*kernel[3]+tmp[4419]*kernel[4]+tmp[4420]*kernel[5]+tmp[4518]*kernel[6]+tmp[4519]*kernel[7]+tmp[4520]*kernel[8];
				ans[4420]<=tmp[4319]*kernel[0]+tmp[4320]*kernel[1]+tmp[4321]*kernel[2]+tmp[4419]*kernel[3]+tmp[4420]*kernel[4]+tmp[4421]*kernel[5]+tmp[4519]*kernel[6]+tmp[4520]*kernel[7]+tmp[4521]*kernel[8];
				ans[4421]<=tmp[4320]*kernel[0]+tmp[4321]*kernel[1]+tmp[4322]*kernel[2]+tmp[4420]*kernel[3]+tmp[4421]*kernel[4]+tmp[4422]*kernel[5]+tmp[4520]*kernel[6]+tmp[4521]*kernel[7]+tmp[4522]*kernel[8];
				ans[4422]<=tmp[4321]*kernel[0]+tmp[4322]*kernel[1]+tmp[4323]*kernel[2]+tmp[4421]*kernel[3]+tmp[4422]*kernel[4]+tmp[4423]*kernel[5]+tmp[4521]*kernel[6]+tmp[4522]*kernel[7]+tmp[4523]*kernel[8];
				ans[4423]<=tmp[4322]*kernel[0]+tmp[4323]*kernel[1]+tmp[4324]*kernel[2]+tmp[4422]*kernel[3]+tmp[4423]*kernel[4]+tmp[4424]*kernel[5]+tmp[4522]*kernel[6]+tmp[4523]*kernel[7]+tmp[4524]*kernel[8];
				ans[4424]<=tmp[4323]*kernel[0]+tmp[4324]*kernel[1]+tmp[4325]*kernel[2]+tmp[4423]*kernel[3]+tmp[4424]*kernel[4]+tmp[4425]*kernel[5]+tmp[4523]*kernel[6]+tmp[4524]*kernel[7]+tmp[4525]*kernel[8];
				ans[4425]<=tmp[4324]*kernel[0]+tmp[4325]*kernel[1]+tmp[4326]*kernel[2]+tmp[4424]*kernel[3]+tmp[4425]*kernel[4]+tmp[4426]*kernel[5]+tmp[4524]*kernel[6]+tmp[4525]*kernel[7]+tmp[4526]*kernel[8];
				ans[4426]<=tmp[4325]*kernel[0]+tmp[4326]*kernel[1]+tmp[4327]*kernel[2]+tmp[4425]*kernel[3]+tmp[4426]*kernel[4]+tmp[4427]*kernel[5]+tmp[4525]*kernel[6]+tmp[4526]*kernel[7]+tmp[4527]*kernel[8];
				ans[4427]<=tmp[4326]*kernel[0]+tmp[4327]*kernel[1]+tmp[4328]*kernel[2]+tmp[4426]*kernel[3]+tmp[4427]*kernel[4]+tmp[4428]*kernel[5]+tmp[4526]*kernel[6]+tmp[4527]*kernel[7]+tmp[4528]*kernel[8];
				ans[4428]<=tmp[4327]*kernel[0]+tmp[4328]*kernel[1]+tmp[4329]*kernel[2]+tmp[4427]*kernel[3]+tmp[4428]*kernel[4]+tmp[4429]*kernel[5]+tmp[4527]*kernel[6]+tmp[4528]*kernel[7]+tmp[4529]*kernel[8];
				ans[4429]<=tmp[4328]*kernel[0]+tmp[4329]*kernel[1]+tmp[4330]*kernel[2]+tmp[4428]*kernel[3]+tmp[4429]*kernel[4]+tmp[4430]*kernel[5]+tmp[4528]*kernel[6]+tmp[4529]*kernel[7]+tmp[4530]*kernel[8];
				ans[4430]<=tmp[4329]*kernel[0]+tmp[4330]*kernel[1]+tmp[4331]*kernel[2]+tmp[4429]*kernel[3]+tmp[4430]*kernel[4]+tmp[4431]*kernel[5]+tmp[4529]*kernel[6]+tmp[4530]*kernel[7]+tmp[4531]*kernel[8];
				ans[4431]<=tmp[4330]*kernel[0]+tmp[4331]*kernel[1]+tmp[4332]*kernel[2]+tmp[4430]*kernel[3]+tmp[4431]*kernel[4]+tmp[4432]*kernel[5]+tmp[4530]*kernel[6]+tmp[4531]*kernel[7]+tmp[4532]*kernel[8];
				ans[4432]<=tmp[4331]*kernel[0]+tmp[4332]*kernel[1]+tmp[4333]*kernel[2]+tmp[4431]*kernel[3]+tmp[4432]*kernel[4]+tmp[4433]*kernel[5]+tmp[4531]*kernel[6]+tmp[4532]*kernel[7]+tmp[4533]*kernel[8];
				ans[4433]<=tmp[4332]*kernel[0]+tmp[4333]*kernel[1]+tmp[4334]*kernel[2]+tmp[4432]*kernel[3]+tmp[4433]*kernel[4]+tmp[4434]*kernel[5]+tmp[4532]*kernel[6]+tmp[4533]*kernel[7]+tmp[4534]*kernel[8];
				ans[4434]<=tmp[4333]*kernel[0]+tmp[4334]*kernel[1]+tmp[4335]*kernel[2]+tmp[4433]*kernel[3]+tmp[4434]*kernel[4]+tmp[4435]*kernel[5]+tmp[4533]*kernel[6]+tmp[4534]*kernel[7]+tmp[4535]*kernel[8];
				ans[4435]<=tmp[4334]*kernel[0]+tmp[4335]*kernel[1]+tmp[4336]*kernel[2]+tmp[4434]*kernel[3]+tmp[4435]*kernel[4]+tmp[4436]*kernel[5]+tmp[4534]*kernel[6]+tmp[4535]*kernel[7]+tmp[4536]*kernel[8];
				ans[4436]<=tmp[4335]*kernel[0]+tmp[4336]*kernel[1]+tmp[4337]*kernel[2]+tmp[4435]*kernel[3]+tmp[4436]*kernel[4]+tmp[4437]*kernel[5]+tmp[4535]*kernel[6]+tmp[4536]*kernel[7]+tmp[4537]*kernel[8];
				ans[4437]<=tmp[4336]*kernel[0]+tmp[4337]*kernel[1]+tmp[4338]*kernel[2]+tmp[4436]*kernel[3]+tmp[4437]*kernel[4]+tmp[4438]*kernel[5]+tmp[4536]*kernel[6]+tmp[4537]*kernel[7]+tmp[4538]*kernel[8];
				ans[4438]<=tmp[4337]*kernel[0]+tmp[4338]*kernel[1]+tmp[4339]*kernel[2]+tmp[4437]*kernel[3]+tmp[4438]*kernel[4]+tmp[4439]*kernel[5]+tmp[4537]*kernel[6]+tmp[4538]*kernel[7]+tmp[4539]*kernel[8];
				ans[4439]<=tmp[4338]*kernel[0]+tmp[4339]*kernel[1]+tmp[4340]*kernel[2]+tmp[4438]*kernel[3]+tmp[4439]*kernel[4]+tmp[4440]*kernel[5]+tmp[4538]*kernel[6]+tmp[4539]*kernel[7]+tmp[4540]*kernel[8];
				ans[4440]<=tmp[4339]*kernel[0]+tmp[4340]*kernel[1]+tmp[4341]*kernel[2]+tmp[4439]*kernel[3]+tmp[4440]*kernel[4]+tmp[4441]*kernel[5]+tmp[4539]*kernel[6]+tmp[4540]*kernel[7]+tmp[4541]*kernel[8];
				ans[4441]<=tmp[4340]*kernel[0]+tmp[4341]*kernel[1]+tmp[4342]*kernel[2]+tmp[4440]*kernel[3]+tmp[4441]*kernel[4]+tmp[4442]*kernel[5]+tmp[4540]*kernel[6]+tmp[4541]*kernel[7]+tmp[4542]*kernel[8];
				ans[4442]<=tmp[4341]*kernel[0]+tmp[4342]*kernel[1]+tmp[4343]*kernel[2]+tmp[4441]*kernel[3]+tmp[4442]*kernel[4]+tmp[4443]*kernel[5]+tmp[4541]*kernel[6]+tmp[4542]*kernel[7]+tmp[4543]*kernel[8];
				ans[4443]<=tmp[4342]*kernel[0]+tmp[4343]*kernel[1]+tmp[4344]*kernel[2]+tmp[4442]*kernel[3]+tmp[4443]*kernel[4]+tmp[4444]*kernel[5]+tmp[4542]*kernel[6]+tmp[4543]*kernel[7]+tmp[4544]*kernel[8];
				ans[4444]<=tmp[4343]*kernel[0]+tmp[4344]*kernel[1]+tmp[4345]*kernel[2]+tmp[4443]*kernel[3]+tmp[4444]*kernel[4]+tmp[4445]*kernel[5]+tmp[4543]*kernel[6]+tmp[4544]*kernel[7]+tmp[4545]*kernel[8];
				ans[4445]<=tmp[4344]*kernel[0]+tmp[4345]*kernel[1]+tmp[4346]*kernel[2]+tmp[4444]*kernel[3]+tmp[4445]*kernel[4]+tmp[4446]*kernel[5]+tmp[4544]*kernel[6]+tmp[4545]*kernel[7]+tmp[4546]*kernel[8];
				ans[4446]<=tmp[4345]*kernel[0]+tmp[4346]*kernel[1]+tmp[4347]*kernel[2]+tmp[4445]*kernel[3]+tmp[4446]*kernel[4]+tmp[4447]*kernel[5]+tmp[4545]*kernel[6]+tmp[4546]*kernel[7]+tmp[4547]*kernel[8];
				ans[4447]<=tmp[4346]*kernel[0]+tmp[4347]*kernel[1]+tmp[4348]*kernel[2]+tmp[4446]*kernel[3]+tmp[4447]*kernel[4]+tmp[4448]*kernel[5]+tmp[4546]*kernel[6]+tmp[4547]*kernel[7]+tmp[4548]*kernel[8];
				ans[4448]<=tmp[4347]*kernel[0]+tmp[4348]*kernel[1]+tmp[4349]*kernel[2]+tmp[4447]*kernel[3]+tmp[4448]*kernel[4]+tmp[4449]*kernel[5]+tmp[4547]*kernel[6]+tmp[4548]*kernel[7]+tmp[4549]*kernel[8];
				ans[4449]<=tmp[4348]*kernel[0]+tmp[4349]*kernel[1]+tmp[4350]*kernel[2]+tmp[4448]*kernel[3]+tmp[4449]*kernel[4]+tmp[4450]*kernel[5]+tmp[4548]*kernel[6]+tmp[4549]*kernel[7]+tmp[4550]*kernel[8];
				ans[4450]<=tmp[4349]*kernel[0]+tmp[4350]*kernel[1]+tmp[4351]*kernel[2]+tmp[4449]*kernel[3]+tmp[4450]*kernel[4]+tmp[4451]*kernel[5]+tmp[4549]*kernel[6]+tmp[4550]*kernel[7]+tmp[4551]*kernel[8];
				ans[4451]<=tmp[4350]*kernel[0]+tmp[4351]*kernel[1]+tmp[4352]*kernel[2]+tmp[4450]*kernel[3]+tmp[4451]*kernel[4]+tmp[4452]*kernel[5]+tmp[4550]*kernel[6]+tmp[4551]*kernel[7]+tmp[4552]*kernel[8];
				ans[4452]<=tmp[4351]*kernel[0]+tmp[4352]*kernel[1]+tmp[4353]*kernel[2]+tmp[4451]*kernel[3]+tmp[4452]*kernel[4]+tmp[4453]*kernel[5]+tmp[4551]*kernel[6]+tmp[4552]*kernel[7]+tmp[4553]*kernel[8];
				ans[4453]<=tmp[4352]*kernel[0]+tmp[4353]*kernel[1]+tmp[4354]*kernel[2]+tmp[4452]*kernel[3]+tmp[4453]*kernel[4]+tmp[4454]*kernel[5]+tmp[4552]*kernel[6]+tmp[4553]*kernel[7]+tmp[4554]*kernel[8];
				ans[4454]<=tmp[4353]*kernel[0]+tmp[4354]*kernel[1]+tmp[4355]*kernel[2]+tmp[4453]*kernel[3]+tmp[4454]*kernel[4]+tmp[4455]*kernel[5]+tmp[4553]*kernel[6]+tmp[4554]*kernel[7]+tmp[4555]*kernel[8];
				ans[4455]<=tmp[4354]*kernel[0]+tmp[4355]*kernel[1]+tmp[4356]*kernel[2]+tmp[4454]*kernel[3]+tmp[4455]*kernel[4]+tmp[4456]*kernel[5]+tmp[4554]*kernel[6]+tmp[4555]*kernel[7]+tmp[4556]*kernel[8];
				ans[4456]<=tmp[4355]*kernel[0]+tmp[4356]*kernel[1]+tmp[4357]*kernel[2]+tmp[4455]*kernel[3]+tmp[4456]*kernel[4]+tmp[4457]*kernel[5]+tmp[4555]*kernel[6]+tmp[4556]*kernel[7]+tmp[4557]*kernel[8];
				ans[4457]<=tmp[4356]*kernel[0]+tmp[4357]*kernel[1]+tmp[4358]*kernel[2]+tmp[4456]*kernel[3]+tmp[4457]*kernel[4]+tmp[4458]*kernel[5]+tmp[4556]*kernel[6]+tmp[4557]*kernel[7]+tmp[4558]*kernel[8];
				ans[4458]<=tmp[4357]*kernel[0]+tmp[4358]*kernel[1]+tmp[4359]*kernel[2]+tmp[4457]*kernel[3]+tmp[4458]*kernel[4]+tmp[4459]*kernel[5]+tmp[4557]*kernel[6]+tmp[4558]*kernel[7]+tmp[4559]*kernel[8];
				ans[4459]<=tmp[4358]*kernel[0]+tmp[4359]*kernel[1]+tmp[4360]*kernel[2]+tmp[4458]*kernel[3]+tmp[4459]*kernel[4]+tmp[4460]*kernel[5]+tmp[4558]*kernel[6]+tmp[4559]*kernel[7]+tmp[4560]*kernel[8];
				ans[4460]<=tmp[4359]*kernel[0]+tmp[4360]*kernel[1]+tmp[4361]*kernel[2]+tmp[4459]*kernel[3]+tmp[4460]*kernel[4]+tmp[4461]*kernel[5]+tmp[4559]*kernel[6]+tmp[4560]*kernel[7]+tmp[4561]*kernel[8];
				ans[4461]<=tmp[4360]*kernel[0]+tmp[4361]*kernel[1]+tmp[4362]*kernel[2]+tmp[4460]*kernel[3]+tmp[4461]*kernel[4]+tmp[4462]*kernel[5]+tmp[4560]*kernel[6]+tmp[4561]*kernel[7]+tmp[4562]*kernel[8];
				ans[4462]<=tmp[4361]*kernel[0]+tmp[4362]*kernel[1]+tmp[4363]*kernel[2]+tmp[4461]*kernel[3]+tmp[4462]*kernel[4]+tmp[4463]*kernel[5]+tmp[4561]*kernel[6]+tmp[4562]*kernel[7]+tmp[4563]*kernel[8];
				ans[4463]<=tmp[4362]*kernel[0]+tmp[4363]*kernel[1]+tmp[4364]*kernel[2]+tmp[4462]*kernel[3]+tmp[4463]*kernel[4]+tmp[4464]*kernel[5]+tmp[4562]*kernel[6]+tmp[4563]*kernel[7]+tmp[4564]*kernel[8];
				ans[4464]<=tmp[4363]*kernel[0]+tmp[4364]*kernel[1]+tmp[4365]*kernel[2]+tmp[4463]*kernel[3]+tmp[4464]*kernel[4]+tmp[4465]*kernel[5]+tmp[4563]*kernel[6]+tmp[4564]*kernel[7]+tmp[4565]*kernel[8];
				ans[4465]<=tmp[4364]*kernel[0]+tmp[4365]*kernel[1]+tmp[4366]*kernel[2]+tmp[4464]*kernel[3]+tmp[4465]*kernel[4]+tmp[4466]*kernel[5]+tmp[4564]*kernel[6]+tmp[4565]*kernel[7]+tmp[4566]*kernel[8];
				ans[4466]<=tmp[4365]*kernel[0]+tmp[4366]*kernel[1]+tmp[4367]*kernel[2]+tmp[4465]*kernel[3]+tmp[4466]*kernel[4]+tmp[4467]*kernel[5]+tmp[4565]*kernel[6]+tmp[4566]*kernel[7]+tmp[4567]*kernel[8];
				ans[4467]<=tmp[4366]*kernel[0]+tmp[4367]*kernel[1]+tmp[4368]*kernel[2]+tmp[4466]*kernel[3]+tmp[4467]*kernel[4]+tmp[4468]*kernel[5]+tmp[4566]*kernel[6]+tmp[4567]*kernel[7]+tmp[4568]*kernel[8];
				ans[4468]<=tmp[4367]*kernel[0]+tmp[4368]*kernel[1]+tmp[4369]*kernel[2]+tmp[4467]*kernel[3]+tmp[4468]*kernel[4]+tmp[4469]*kernel[5]+tmp[4567]*kernel[6]+tmp[4568]*kernel[7]+tmp[4569]*kernel[8];
				ans[4469]<=tmp[4368]*kernel[0]+tmp[4369]*kernel[1]+tmp[4370]*kernel[2]+tmp[4468]*kernel[3]+tmp[4469]*kernel[4]+tmp[4470]*kernel[5]+tmp[4568]*kernel[6]+tmp[4569]*kernel[7]+tmp[4570]*kernel[8];
				ans[4470]<=tmp[4369]*kernel[0]+tmp[4370]*kernel[1]+tmp[4371]*kernel[2]+tmp[4469]*kernel[3]+tmp[4470]*kernel[4]+tmp[4471]*kernel[5]+tmp[4569]*kernel[6]+tmp[4570]*kernel[7]+tmp[4571]*kernel[8];
				ans[4471]<=tmp[4370]*kernel[0]+tmp[4371]*kernel[1]+tmp[4372]*kernel[2]+tmp[4470]*kernel[3]+tmp[4471]*kernel[4]+tmp[4472]*kernel[5]+tmp[4570]*kernel[6]+tmp[4571]*kernel[7]+tmp[4572]*kernel[8];
				ans[4472]<=tmp[4371]*kernel[0]+tmp[4372]*kernel[1]+tmp[4373]*kernel[2]+tmp[4471]*kernel[3]+tmp[4472]*kernel[4]+tmp[4473]*kernel[5]+tmp[4571]*kernel[6]+tmp[4572]*kernel[7]+tmp[4573]*kernel[8];
				ans[4473]<=tmp[4372]*kernel[0]+tmp[4373]*kernel[1]+tmp[4374]*kernel[2]+tmp[4472]*kernel[3]+tmp[4473]*kernel[4]+tmp[4474]*kernel[5]+tmp[4572]*kernel[6]+tmp[4573]*kernel[7]+tmp[4574]*kernel[8];
				ans[4474]<=tmp[4373]*kernel[0]+tmp[4374]*kernel[1]+tmp[4375]*kernel[2]+tmp[4473]*kernel[3]+tmp[4474]*kernel[4]+tmp[4475]*kernel[5]+tmp[4573]*kernel[6]+tmp[4574]*kernel[7]+tmp[4575]*kernel[8];
				ans[4475]<=tmp[4374]*kernel[0]+tmp[4375]*kernel[1]+tmp[4376]*kernel[2]+tmp[4474]*kernel[3]+tmp[4475]*kernel[4]+tmp[4476]*kernel[5]+tmp[4574]*kernel[6]+tmp[4575]*kernel[7]+tmp[4576]*kernel[8];
				ans[4476]<=tmp[4375]*kernel[0]+tmp[4376]*kernel[1]+tmp[4377]*kernel[2]+tmp[4475]*kernel[3]+tmp[4476]*kernel[4]+tmp[4477]*kernel[5]+tmp[4575]*kernel[6]+tmp[4576]*kernel[7]+tmp[4577]*kernel[8];
				ans[4477]<=tmp[4376]*kernel[0]+tmp[4377]*kernel[1]+tmp[4378]*kernel[2]+tmp[4476]*kernel[3]+tmp[4477]*kernel[4]+tmp[4478]*kernel[5]+tmp[4576]*kernel[6]+tmp[4577]*kernel[7]+tmp[4578]*kernel[8];
				ans[4478]<=tmp[4377]*kernel[0]+tmp[4378]*kernel[1]+tmp[4379]*kernel[2]+tmp[4477]*kernel[3]+tmp[4478]*kernel[4]+tmp[4479]*kernel[5]+tmp[4577]*kernel[6]+tmp[4578]*kernel[7]+tmp[4579]*kernel[8];
				ans[4479]<=tmp[4378]*kernel[0]+tmp[4379]*kernel[1]+tmp[4380]*kernel[2]+tmp[4478]*kernel[3]+tmp[4479]*kernel[4]+tmp[4480]*kernel[5]+tmp[4578]*kernel[6]+tmp[4579]*kernel[7]+tmp[4580]*kernel[8];
				ans[4480]<=tmp[4379]*kernel[0]+tmp[4380]*kernel[1]+tmp[4381]*kernel[2]+tmp[4479]*kernel[3]+tmp[4480]*kernel[4]+tmp[4481]*kernel[5]+tmp[4579]*kernel[6]+tmp[4580]*kernel[7]+tmp[4581]*kernel[8];
				ans[4481]<=tmp[4380]*kernel[0]+tmp[4381]*kernel[1]+tmp[4382]*kernel[2]+tmp[4480]*kernel[3]+tmp[4481]*kernel[4]+tmp[4482]*kernel[5]+tmp[4580]*kernel[6]+tmp[4581]*kernel[7]+tmp[4582]*kernel[8];
				ans[4482]<=tmp[4381]*kernel[0]+tmp[4382]*kernel[1]+tmp[4383]*kernel[2]+tmp[4481]*kernel[3]+tmp[4482]*kernel[4]+tmp[4483]*kernel[5]+tmp[4581]*kernel[6]+tmp[4582]*kernel[7]+tmp[4583]*kernel[8];
				ans[4483]<=tmp[4382]*kernel[0]+tmp[4383]*kernel[1]+tmp[4384]*kernel[2]+tmp[4482]*kernel[3]+tmp[4483]*kernel[4]+tmp[4484]*kernel[5]+tmp[4582]*kernel[6]+tmp[4583]*kernel[7]+tmp[4584]*kernel[8];
				ans[4484]<=tmp[4383]*kernel[0]+tmp[4384]*kernel[1]+tmp[4385]*kernel[2]+tmp[4483]*kernel[3]+tmp[4484]*kernel[4]+tmp[4485]*kernel[5]+tmp[4583]*kernel[6]+tmp[4584]*kernel[7]+tmp[4585]*kernel[8];
				ans[4485]<=tmp[4384]*kernel[0]+tmp[4385]*kernel[1]+tmp[4386]*kernel[2]+tmp[4484]*kernel[3]+tmp[4485]*kernel[4]+tmp[4486]*kernel[5]+tmp[4584]*kernel[6]+tmp[4585]*kernel[7]+tmp[4586]*kernel[8];
				ans[4486]<=tmp[4385]*kernel[0]+tmp[4386]*kernel[1]+tmp[4387]*kernel[2]+tmp[4485]*kernel[3]+tmp[4486]*kernel[4]+tmp[4487]*kernel[5]+tmp[4585]*kernel[6]+tmp[4586]*kernel[7]+tmp[4587]*kernel[8];
				ans[4487]<=tmp[4386]*kernel[0]+tmp[4387]*kernel[1]+tmp[4388]*kernel[2]+tmp[4486]*kernel[3]+tmp[4487]*kernel[4]+tmp[4488]*kernel[5]+tmp[4586]*kernel[6]+tmp[4587]*kernel[7]+tmp[4588]*kernel[8];
				ans[4488]<=tmp[4387]*kernel[0]+tmp[4388]*kernel[1]+tmp[4389]*kernel[2]+tmp[4487]*kernel[3]+tmp[4488]*kernel[4]+tmp[4489]*kernel[5]+tmp[4587]*kernel[6]+tmp[4588]*kernel[7]+tmp[4589]*kernel[8];
				ans[4489]<=tmp[4388]*kernel[0]+tmp[4389]*kernel[1]+tmp[4390]*kernel[2]+tmp[4488]*kernel[3]+tmp[4489]*kernel[4]+tmp[4490]*kernel[5]+tmp[4588]*kernel[6]+tmp[4589]*kernel[7]+tmp[4590]*kernel[8];
				ans[4490]<=tmp[4389]*kernel[0]+tmp[4390]*kernel[1]+tmp[4391]*kernel[2]+tmp[4489]*kernel[3]+tmp[4490]*kernel[4]+tmp[4491]*kernel[5]+tmp[4589]*kernel[6]+tmp[4590]*kernel[7]+tmp[4591]*kernel[8];
				ans[4491]<=tmp[4390]*kernel[0]+tmp[4391]*kernel[1]+tmp[4392]*kernel[2]+tmp[4490]*kernel[3]+tmp[4491]*kernel[4]+tmp[4492]*kernel[5]+tmp[4590]*kernel[6]+tmp[4591]*kernel[7]+tmp[4592]*kernel[8];
				ans[4492]<=tmp[4391]*kernel[0]+tmp[4392]*kernel[1]+tmp[4393]*kernel[2]+tmp[4491]*kernel[3]+tmp[4492]*kernel[4]+tmp[4493]*kernel[5]+tmp[4591]*kernel[6]+tmp[4592]*kernel[7]+tmp[4593]*kernel[8];
				ans[4493]<=tmp[4392]*kernel[0]+tmp[4393]*kernel[1]+tmp[4394]*kernel[2]+tmp[4492]*kernel[3]+tmp[4493]*kernel[4]+tmp[4494]*kernel[5]+tmp[4592]*kernel[6]+tmp[4593]*kernel[7]+tmp[4594]*kernel[8];
				ans[4494]<=tmp[4393]*kernel[0]+tmp[4394]*kernel[1]+tmp[4395]*kernel[2]+tmp[4493]*kernel[3]+tmp[4494]*kernel[4]+tmp[4495]*kernel[5]+tmp[4593]*kernel[6]+tmp[4594]*kernel[7]+tmp[4595]*kernel[8];
				ans[4495]<=tmp[4394]*kernel[0]+tmp[4395]*kernel[1]+tmp[4396]*kernel[2]+tmp[4494]*kernel[3]+tmp[4495]*kernel[4]+tmp[4496]*kernel[5]+tmp[4594]*kernel[6]+tmp[4595]*kernel[7]+tmp[4596]*kernel[8];
				ans[4496]<=tmp[4395]*kernel[0]+tmp[4396]*kernel[1]+tmp[4397]*kernel[2]+tmp[4495]*kernel[3]+tmp[4496]*kernel[4]+tmp[4497]*kernel[5]+tmp[4595]*kernel[6]+tmp[4596]*kernel[7]+tmp[4597]*kernel[8];
				ans[4497]<=tmp[4396]*kernel[0]+tmp[4397]*kernel[1]+tmp[4398]*kernel[2]+tmp[4496]*kernel[3]+tmp[4497]*kernel[4]+tmp[4498]*kernel[5]+tmp[4596]*kernel[6]+tmp[4597]*kernel[7]+tmp[4598]*kernel[8];
				ans[4498]<=tmp[4397]*kernel[0]+tmp[4398]*kernel[1]+tmp[4399]*kernel[2]+tmp[4497]*kernel[3]+tmp[4498]*kernel[4]+tmp[4499]*kernel[5]+tmp[4597]*kernel[6]+tmp[4598]*kernel[7]+tmp[4599]*kernel[8];
				ans[4499]<=tmp[4398]*kernel[0]+tmp[4399]*kernel[1]+tmp[4498]*kernel[3]+tmp[4499]*kernel[4]+tmp[4598]*kernel[6]+tmp[4599]*kernel[7];
				ans[4500]<=tmp[4400]*kernel[1]+tmp[4401]*kernel[2]+tmp[4500]*kernel[4]+tmp[4501]*kernel[5]+tmp[4600]*kernel[7]+tmp[4601]*kernel[8];
				ans[4501]<=tmp[4400]*kernel[0]+tmp[4401]*kernel[1]+tmp[4402]*kernel[2]+tmp[4500]*kernel[3]+tmp[4501]*kernel[4]+tmp[4502]*kernel[5]+tmp[4600]*kernel[6]+tmp[4601]*kernel[7]+tmp[4602]*kernel[8];
				ans[4502]<=tmp[4401]*kernel[0]+tmp[4402]*kernel[1]+tmp[4403]*kernel[2]+tmp[4501]*kernel[3]+tmp[4502]*kernel[4]+tmp[4503]*kernel[5]+tmp[4601]*kernel[6]+tmp[4602]*kernel[7]+tmp[4603]*kernel[8];
				ans[4503]<=tmp[4402]*kernel[0]+tmp[4403]*kernel[1]+tmp[4404]*kernel[2]+tmp[4502]*kernel[3]+tmp[4503]*kernel[4]+tmp[4504]*kernel[5]+tmp[4602]*kernel[6]+tmp[4603]*kernel[7]+tmp[4604]*kernel[8];
				ans[4504]<=tmp[4403]*kernel[0]+tmp[4404]*kernel[1]+tmp[4405]*kernel[2]+tmp[4503]*kernel[3]+tmp[4504]*kernel[4]+tmp[4505]*kernel[5]+tmp[4603]*kernel[6]+tmp[4604]*kernel[7]+tmp[4605]*kernel[8];
				ans[4505]<=tmp[4404]*kernel[0]+tmp[4405]*kernel[1]+tmp[4406]*kernel[2]+tmp[4504]*kernel[3]+tmp[4505]*kernel[4]+tmp[4506]*kernel[5]+tmp[4604]*kernel[6]+tmp[4605]*kernel[7]+tmp[4606]*kernel[8];
				ans[4506]<=tmp[4405]*kernel[0]+tmp[4406]*kernel[1]+tmp[4407]*kernel[2]+tmp[4505]*kernel[3]+tmp[4506]*kernel[4]+tmp[4507]*kernel[5]+tmp[4605]*kernel[6]+tmp[4606]*kernel[7]+tmp[4607]*kernel[8];
				ans[4507]<=tmp[4406]*kernel[0]+tmp[4407]*kernel[1]+tmp[4408]*kernel[2]+tmp[4506]*kernel[3]+tmp[4507]*kernel[4]+tmp[4508]*kernel[5]+tmp[4606]*kernel[6]+tmp[4607]*kernel[7]+tmp[4608]*kernel[8];
				ans[4508]<=tmp[4407]*kernel[0]+tmp[4408]*kernel[1]+tmp[4409]*kernel[2]+tmp[4507]*kernel[3]+tmp[4508]*kernel[4]+tmp[4509]*kernel[5]+tmp[4607]*kernel[6]+tmp[4608]*kernel[7]+tmp[4609]*kernel[8];
				ans[4509]<=tmp[4408]*kernel[0]+tmp[4409]*kernel[1]+tmp[4410]*kernel[2]+tmp[4508]*kernel[3]+tmp[4509]*kernel[4]+tmp[4510]*kernel[5]+tmp[4608]*kernel[6]+tmp[4609]*kernel[7]+tmp[4610]*kernel[8];
				ans[4510]<=tmp[4409]*kernel[0]+tmp[4410]*kernel[1]+tmp[4411]*kernel[2]+tmp[4509]*kernel[3]+tmp[4510]*kernel[4]+tmp[4511]*kernel[5]+tmp[4609]*kernel[6]+tmp[4610]*kernel[7]+tmp[4611]*kernel[8];
				ans[4511]<=tmp[4410]*kernel[0]+tmp[4411]*kernel[1]+tmp[4412]*kernel[2]+tmp[4510]*kernel[3]+tmp[4511]*kernel[4]+tmp[4512]*kernel[5]+tmp[4610]*kernel[6]+tmp[4611]*kernel[7]+tmp[4612]*kernel[8];
				ans[4512]<=tmp[4411]*kernel[0]+tmp[4412]*kernel[1]+tmp[4413]*kernel[2]+tmp[4511]*kernel[3]+tmp[4512]*kernel[4]+tmp[4513]*kernel[5]+tmp[4611]*kernel[6]+tmp[4612]*kernel[7]+tmp[4613]*kernel[8];
				ans[4513]<=tmp[4412]*kernel[0]+tmp[4413]*kernel[1]+tmp[4414]*kernel[2]+tmp[4512]*kernel[3]+tmp[4513]*kernel[4]+tmp[4514]*kernel[5]+tmp[4612]*kernel[6]+tmp[4613]*kernel[7]+tmp[4614]*kernel[8];
				ans[4514]<=tmp[4413]*kernel[0]+tmp[4414]*kernel[1]+tmp[4415]*kernel[2]+tmp[4513]*kernel[3]+tmp[4514]*kernel[4]+tmp[4515]*kernel[5]+tmp[4613]*kernel[6]+tmp[4614]*kernel[7]+tmp[4615]*kernel[8];
				ans[4515]<=tmp[4414]*kernel[0]+tmp[4415]*kernel[1]+tmp[4416]*kernel[2]+tmp[4514]*kernel[3]+tmp[4515]*kernel[4]+tmp[4516]*kernel[5]+tmp[4614]*kernel[6]+tmp[4615]*kernel[7]+tmp[4616]*kernel[8];
				ans[4516]<=tmp[4415]*kernel[0]+tmp[4416]*kernel[1]+tmp[4417]*kernel[2]+tmp[4515]*kernel[3]+tmp[4516]*kernel[4]+tmp[4517]*kernel[5]+tmp[4615]*kernel[6]+tmp[4616]*kernel[7]+tmp[4617]*kernel[8];
				ans[4517]<=tmp[4416]*kernel[0]+tmp[4417]*kernel[1]+tmp[4418]*kernel[2]+tmp[4516]*kernel[3]+tmp[4517]*kernel[4]+tmp[4518]*kernel[5]+tmp[4616]*kernel[6]+tmp[4617]*kernel[7]+tmp[4618]*kernel[8];
				ans[4518]<=tmp[4417]*kernel[0]+tmp[4418]*kernel[1]+tmp[4419]*kernel[2]+tmp[4517]*kernel[3]+tmp[4518]*kernel[4]+tmp[4519]*kernel[5]+tmp[4617]*kernel[6]+tmp[4618]*kernel[7]+tmp[4619]*kernel[8];
				ans[4519]<=tmp[4418]*kernel[0]+tmp[4419]*kernel[1]+tmp[4420]*kernel[2]+tmp[4518]*kernel[3]+tmp[4519]*kernel[4]+tmp[4520]*kernel[5]+tmp[4618]*kernel[6]+tmp[4619]*kernel[7]+tmp[4620]*kernel[8];
				ans[4520]<=tmp[4419]*kernel[0]+tmp[4420]*kernel[1]+tmp[4421]*kernel[2]+tmp[4519]*kernel[3]+tmp[4520]*kernel[4]+tmp[4521]*kernel[5]+tmp[4619]*kernel[6]+tmp[4620]*kernel[7]+tmp[4621]*kernel[8];
				ans[4521]<=tmp[4420]*kernel[0]+tmp[4421]*kernel[1]+tmp[4422]*kernel[2]+tmp[4520]*kernel[3]+tmp[4521]*kernel[4]+tmp[4522]*kernel[5]+tmp[4620]*kernel[6]+tmp[4621]*kernel[7]+tmp[4622]*kernel[8];
				ans[4522]<=tmp[4421]*kernel[0]+tmp[4422]*kernel[1]+tmp[4423]*kernel[2]+tmp[4521]*kernel[3]+tmp[4522]*kernel[4]+tmp[4523]*kernel[5]+tmp[4621]*kernel[6]+tmp[4622]*kernel[7]+tmp[4623]*kernel[8];
				ans[4523]<=tmp[4422]*kernel[0]+tmp[4423]*kernel[1]+tmp[4424]*kernel[2]+tmp[4522]*kernel[3]+tmp[4523]*kernel[4]+tmp[4524]*kernel[5]+tmp[4622]*kernel[6]+tmp[4623]*kernel[7]+tmp[4624]*kernel[8];
				ans[4524]<=tmp[4423]*kernel[0]+tmp[4424]*kernel[1]+tmp[4425]*kernel[2]+tmp[4523]*kernel[3]+tmp[4524]*kernel[4]+tmp[4525]*kernel[5]+tmp[4623]*kernel[6]+tmp[4624]*kernel[7]+tmp[4625]*kernel[8];
				ans[4525]<=tmp[4424]*kernel[0]+tmp[4425]*kernel[1]+tmp[4426]*kernel[2]+tmp[4524]*kernel[3]+tmp[4525]*kernel[4]+tmp[4526]*kernel[5]+tmp[4624]*kernel[6]+tmp[4625]*kernel[7]+tmp[4626]*kernel[8];
				ans[4526]<=tmp[4425]*kernel[0]+tmp[4426]*kernel[1]+tmp[4427]*kernel[2]+tmp[4525]*kernel[3]+tmp[4526]*kernel[4]+tmp[4527]*kernel[5]+tmp[4625]*kernel[6]+tmp[4626]*kernel[7]+tmp[4627]*kernel[8];
				ans[4527]<=tmp[4426]*kernel[0]+tmp[4427]*kernel[1]+tmp[4428]*kernel[2]+tmp[4526]*kernel[3]+tmp[4527]*kernel[4]+tmp[4528]*kernel[5]+tmp[4626]*kernel[6]+tmp[4627]*kernel[7]+tmp[4628]*kernel[8];
				ans[4528]<=tmp[4427]*kernel[0]+tmp[4428]*kernel[1]+tmp[4429]*kernel[2]+tmp[4527]*kernel[3]+tmp[4528]*kernel[4]+tmp[4529]*kernel[5]+tmp[4627]*kernel[6]+tmp[4628]*kernel[7]+tmp[4629]*kernel[8];
				ans[4529]<=tmp[4428]*kernel[0]+tmp[4429]*kernel[1]+tmp[4430]*kernel[2]+tmp[4528]*kernel[3]+tmp[4529]*kernel[4]+tmp[4530]*kernel[5]+tmp[4628]*kernel[6]+tmp[4629]*kernel[7]+tmp[4630]*kernel[8];
				ans[4530]<=tmp[4429]*kernel[0]+tmp[4430]*kernel[1]+tmp[4431]*kernel[2]+tmp[4529]*kernel[3]+tmp[4530]*kernel[4]+tmp[4531]*kernel[5]+tmp[4629]*kernel[6]+tmp[4630]*kernel[7]+tmp[4631]*kernel[8];
				ans[4531]<=tmp[4430]*kernel[0]+tmp[4431]*kernel[1]+tmp[4432]*kernel[2]+tmp[4530]*kernel[3]+tmp[4531]*kernel[4]+tmp[4532]*kernel[5]+tmp[4630]*kernel[6]+tmp[4631]*kernel[7]+tmp[4632]*kernel[8];
				ans[4532]<=tmp[4431]*kernel[0]+tmp[4432]*kernel[1]+tmp[4433]*kernel[2]+tmp[4531]*kernel[3]+tmp[4532]*kernel[4]+tmp[4533]*kernel[5]+tmp[4631]*kernel[6]+tmp[4632]*kernel[7]+tmp[4633]*kernel[8];
				ans[4533]<=tmp[4432]*kernel[0]+tmp[4433]*kernel[1]+tmp[4434]*kernel[2]+tmp[4532]*kernel[3]+tmp[4533]*kernel[4]+tmp[4534]*kernel[5]+tmp[4632]*kernel[6]+tmp[4633]*kernel[7]+tmp[4634]*kernel[8];
				ans[4534]<=tmp[4433]*kernel[0]+tmp[4434]*kernel[1]+tmp[4435]*kernel[2]+tmp[4533]*kernel[3]+tmp[4534]*kernel[4]+tmp[4535]*kernel[5]+tmp[4633]*kernel[6]+tmp[4634]*kernel[7]+tmp[4635]*kernel[8];
				ans[4535]<=tmp[4434]*kernel[0]+tmp[4435]*kernel[1]+tmp[4436]*kernel[2]+tmp[4534]*kernel[3]+tmp[4535]*kernel[4]+tmp[4536]*kernel[5]+tmp[4634]*kernel[6]+tmp[4635]*kernel[7]+tmp[4636]*kernel[8];
				ans[4536]<=tmp[4435]*kernel[0]+tmp[4436]*kernel[1]+tmp[4437]*kernel[2]+tmp[4535]*kernel[3]+tmp[4536]*kernel[4]+tmp[4537]*kernel[5]+tmp[4635]*kernel[6]+tmp[4636]*kernel[7]+tmp[4637]*kernel[8];
				ans[4537]<=tmp[4436]*kernel[0]+tmp[4437]*kernel[1]+tmp[4438]*kernel[2]+tmp[4536]*kernel[3]+tmp[4537]*kernel[4]+tmp[4538]*kernel[5]+tmp[4636]*kernel[6]+tmp[4637]*kernel[7]+tmp[4638]*kernel[8];
				ans[4538]<=tmp[4437]*kernel[0]+tmp[4438]*kernel[1]+tmp[4439]*kernel[2]+tmp[4537]*kernel[3]+tmp[4538]*kernel[4]+tmp[4539]*kernel[5]+tmp[4637]*kernel[6]+tmp[4638]*kernel[7]+tmp[4639]*kernel[8];
				ans[4539]<=tmp[4438]*kernel[0]+tmp[4439]*kernel[1]+tmp[4440]*kernel[2]+tmp[4538]*kernel[3]+tmp[4539]*kernel[4]+tmp[4540]*kernel[5]+tmp[4638]*kernel[6]+tmp[4639]*kernel[7]+tmp[4640]*kernel[8];
				ans[4540]<=tmp[4439]*kernel[0]+tmp[4440]*kernel[1]+tmp[4441]*kernel[2]+tmp[4539]*kernel[3]+tmp[4540]*kernel[4]+tmp[4541]*kernel[5]+tmp[4639]*kernel[6]+tmp[4640]*kernel[7]+tmp[4641]*kernel[8];
				ans[4541]<=tmp[4440]*kernel[0]+tmp[4441]*kernel[1]+tmp[4442]*kernel[2]+tmp[4540]*kernel[3]+tmp[4541]*kernel[4]+tmp[4542]*kernel[5]+tmp[4640]*kernel[6]+tmp[4641]*kernel[7]+tmp[4642]*kernel[8];
				ans[4542]<=tmp[4441]*kernel[0]+tmp[4442]*kernel[1]+tmp[4443]*kernel[2]+tmp[4541]*kernel[3]+tmp[4542]*kernel[4]+tmp[4543]*kernel[5]+tmp[4641]*kernel[6]+tmp[4642]*kernel[7]+tmp[4643]*kernel[8];
				ans[4543]<=tmp[4442]*kernel[0]+tmp[4443]*kernel[1]+tmp[4444]*kernel[2]+tmp[4542]*kernel[3]+tmp[4543]*kernel[4]+tmp[4544]*kernel[5]+tmp[4642]*kernel[6]+tmp[4643]*kernel[7]+tmp[4644]*kernel[8];
				ans[4544]<=tmp[4443]*kernel[0]+tmp[4444]*kernel[1]+tmp[4445]*kernel[2]+tmp[4543]*kernel[3]+tmp[4544]*kernel[4]+tmp[4545]*kernel[5]+tmp[4643]*kernel[6]+tmp[4644]*kernel[7]+tmp[4645]*kernel[8];
				ans[4545]<=tmp[4444]*kernel[0]+tmp[4445]*kernel[1]+tmp[4446]*kernel[2]+tmp[4544]*kernel[3]+tmp[4545]*kernel[4]+tmp[4546]*kernel[5]+tmp[4644]*kernel[6]+tmp[4645]*kernel[7]+tmp[4646]*kernel[8];
				ans[4546]<=tmp[4445]*kernel[0]+tmp[4446]*kernel[1]+tmp[4447]*kernel[2]+tmp[4545]*kernel[3]+tmp[4546]*kernel[4]+tmp[4547]*kernel[5]+tmp[4645]*kernel[6]+tmp[4646]*kernel[7]+tmp[4647]*kernel[8];
				ans[4547]<=tmp[4446]*kernel[0]+tmp[4447]*kernel[1]+tmp[4448]*kernel[2]+tmp[4546]*kernel[3]+tmp[4547]*kernel[4]+tmp[4548]*kernel[5]+tmp[4646]*kernel[6]+tmp[4647]*kernel[7]+tmp[4648]*kernel[8];
				ans[4548]<=tmp[4447]*kernel[0]+tmp[4448]*kernel[1]+tmp[4449]*kernel[2]+tmp[4547]*kernel[3]+tmp[4548]*kernel[4]+tmp[4549]*kernel[5]+tmp[4647]*kernel[6]+tmp[4648]*kernel[7]+tmp[4649]*kernel[8];
				ans[4549]<=tmp[4448]*kernel[0]+tmp[4449]*kernel[1]+tmp[4450]*kernel[2]+tmp[4548]*kernel[3]+tmp[4549]*kernel[4]+tmp[4550]*kernel[5]+tmp[4648]*kernel[6]+tmp[4649]*kernel[7]+tmp[4650]*kernel[8];
				ans[4550]<=tmp[4449]*kernel[0]+tmp[4450]*kernel[1]+tmp[4451]*kernel[2]+tmp[4549]*kernel[3]+tmp[4550]*kernel[4]+tmp[4551]*kernel[5]+tmp[4649]*kernel[6]+tmp[4650]*kernel[7]+tmp[4651]*kernel[8];
				ans[4551]<=tmp[4450]*kernel[0]+tmp[4451]*kernel[1]+tmp[4452]*kernel[2]+tmp[4550]*kernel[3]+tmp[4551]*kernel[4]+tmp[4552]*kernel[5]+tmp[4650]*kernel[6]+tmp[4651]*kernel[7]+tmp[4652]*kernel[8];
				ans[4552]<=tmp[4451]*kernel[0]+tmp[4452]*kernel[1]+tmp[4453]*kernel[2]+tmp[4551]*kernel[3]+tmp[4552]*kernel[4]+tmp[4553]*kernel[5]+tmp[4651]*kernel[6]+tmp[4652]*kernel[7]+tmp[4653]*kernel[8];
				ans[4553]<=tmp[4452]*kernel[0]+tmp[4453]*kernel[1]+tmp[4454]*kernel[2]+tmp[4552]*kernel[3]+tmp[4553]*kernel[4]+tmp[4554]*kernel[5]+tmp[4652]*kernel[6]+tmp[4653]*kernel[7]+tmp[4654]*kernel[8];
				ans[4554]<=tmp[4453]*kernel[0]+tmp[4454]*kernel[1]+tmp[4455]*kernel[2]+tmp[4553]*kernel[3]+tmp[4554]*kernel[4]+tmp[4555]*kernel[5]+tmp[4653]*kernel[6]+tmp[4654]*kernel[7]+tmp[4655]*kernel[8];
				ans[4555]<=tmp[4454]*kernel[0]+tmp[4455]*kernel[1]+tmp[4456]*kernel[2]+tmp[4554]*kernel[3]+tmp[4555]*kernel[4]+tmp[4556]*kernel[5]+tmp[4654]*kernel[6]+tmp[4655]*kernel[7]+tmp[4656]*kernel[8];
				ans[4556]<=tmp[4455]*kernel[0]+tmp[4456]*kernel[1]+tmp[4457]*kernel[2]+tmp[4555]*kernel[3]+tmp[4556]*kernel[4]+tmp[4557]*kernel[5]+tmp[4655]*kernel[6]+tmp[4656]*kernel[7]+tmp[4657]*kernel[8];
				ans[4557]<=tmp[4456]*kernel[0]+tmp[4457]*kernel[1]+tmp[4458]*kernel[2]+tmp[4556]*kernel[3]+tmp[4557]*kernel[4]+tmp[4558]*kernel[5]+tmp[4656]*kernel[6]+tmp[4657]*kernel[7]+tmp[4658]*kernel[8];
				ans[4558]<=tmp[4457]*kernel[0]+tmp[4458]*kernel[1]+tmp[4459]*kernel[2]+tmp[4557]*kernel[3]+tmp[4558]*kernel[4]+tmp[4559]*kernel[5]+tmp[4657]*kernel[6]+tmp[4658]*kernel[7]+tmp[4659]*kernel[8];
				ans[4559]<=tmp[4458]*kernel[0]+tmp[4459]*kernel[1]+tmp[4460]*kernel[2]+tmp[4558]*kernel[3]+tmp[4559]*kernel[4]+tmp[4560]*kernel[5]+tmp[4658]*kernel[6]+tmp[4659]*kernel[7]+tmp[4660]*kernel[8];
				ans[4560]<=tmp[4459]*kernel[0]+tmp[4460]*kernel[1]+tmp[4461]*kernel[2]+tmp[4559]*kernel[3]+tmp[4560]*kernel[4]+tmp[4561]*kernel[5]+tmp[4659]*kernel[6]+tmp[4660]*kernel[7]+tmp[4661]*kernel[8];
				ans[4561]<=tmp[4460]*kernel[0]+tmp[4461]*kernel[1]+tmp[4462]*kernel[2]+tmp[4560]*kernel[3]+tmp[4561]*kernel[4]+tmp[4562]*kernel[5]+tmp[4660]*kernel[6]+tmp[4661]*kernel[7]+tmp[4662]*kernel[8];
				ans[4562]<=tmp[4461]*kernel[0]+tmp[4462]*kernel[1]+tmp[4463]*kernel[2]+tmp[4561]*kernel[3]+tmp[4562]*kernel[4]+tmp[4563]*kernel[5]+tmp[4661]*kernel[6]+tmp[4662]*kernel[7]+tmp[4663]*kernel[8];
				ans[4563]<=tmp[4462]*kernel[0]+tmp[4463]*kernel[1]+tmp[4464]*kernel[2]+tmp[4562]*kernel[3]+tmp[4563]*kernel[4]+tmp[4564]*kernel[5]+tmp[4662]*kernel[6]+tmp[4663]*kernel[7]+tmp[4664]*kernel[8];
				ans[4564]<=tmp[4463]*kernel[0]+tmp[4464]*kernel[1]+tmp[4465]*kernel[2]+tmp[4563]*kernel[3]+tmp[4564]*kernel[4]+tmp[4565]*kernel[5]+tmp[4663]*kernel[6]+tmp[4664]*kernel[7]+tmp[4665]*kernel[8];
				ans[4565]<=tmp[4464]*kernel[0]+tmp[4465]*kernel[1]+tmp[4466]*kernel[2]+tmp[4564]*kernel[3]+tmp[4565]*kernel[4]+tmp[4566]*kernel[5]+tmp[4664]*kernel[6]+tmp[4665]*kernel[7]+tmp[4666]*kernel[8];
				ans[4566]<=tmp[4465]*kernel[0]+tmp[4466]*kernel[1]+tmp[4467]*kernel[2]+tmp[4565]*kernel[3]+tmp[4566]*kernel[4]+tmp[4567]*kernel[5]+tmp[4665]*kernel[6]+tmp[4666]*kernel[7]+tmp[4667]*kernel[8];
				ans[4567]<=tmp[4466]*kernel[0]+tmp[4467]*kernel[1]+tmp[4468]*kernel[2]+tmp[4566]*kernel[3]+tmp[4567]*kernel[4]+tmp[4568]*kernel[5]+tmp[4666]*kernel[6]+tmp[4667]*kernel[7]+tmp[4668]*kernel[8];
				ans[4568]<=tmp[4467]*kernel[0]+tmp[4468]*kernel[1]+tmp[4469]*kernel[2]+tmp[4567]*kernel[3]+tmp[4568]*kernel[4]+tmp[4569]*kernel[5]+tmp[4667]*kernel[6]+tmp[4668]*kernel[7]+tmp[4669]*kernel[8];
				ans[4569]<=tmp[4468]*kernel[0]+tmp[4469]*kernel[1]+tmp[4470]*kernel[2]+tmp[4568]*kernel[3]+tmp[4569]*kernel[4]+tmp[4570]*kernel[5]+tmp[4668]*kernel[6]+tmp[4669]*kernel[7]+tmp[4670]*kernel[8];
				ans[4570]<=tmp[4469]*kernel[0]+tmp[4470]*kernel[1]+tmp[4471]*kernel[2]+tmp[4569]*kernel[3]+tmp[4570]*kernel[4]+tmp[4571]*kernel[5]+tmp[4669]*kernel[6]+tmp[4670]*kernel[7]+tmp[4671]*kernel[8];
				ans[4571]<=tmp[4470]*kernel[0]+tmp[4471]*kernel[1]+tmp[4472]*kernel[2]+tmp[4570]*kernel[3]+tmp[4571]*kernel[4]+tmp[4572]*kernel[5]+tmp[4670]*kernel[6]+tmp[4671]*kernel[7]+tmp[4672]*kernel[8];
				ans[4572]<=tmp[4471]*kernel[0]+tmp[4472]*kernel[1]+tmp[4473]*kernel[2]+tmp[4571]*kernel[3]+tmp[4572]*kernel[4]+tmp[4573]*kernel[5]+tmp[4671]*kernel[6]+tmp[4672]*kernel[7]+tmp[4673]*kernel[8];
				ans[4573]<=tmp[4472]*kernel[0]+tmp[4473]*kernel[1]+tmp[4474]*kernel[2]+tmp[4572]*kernel[3]+tmp[4573]*kernel[4]+tmp[4574]*kernel[5]+tmp[4672]*kernel[6]+tmp[4673]*kernel[7]+tmp[4674]*kernel[8];
				ans[4574]<=tmp[4473]*kernel[0]+tmp[4474]*kernel[1]+tmp[4475]*kernel[2]+tmp[4573]*kernel[3]+tmp[4574]*kernel[4]+tmp[4575]*kernel[5]+tmp[4673]*kernel[6]+tmp[4674]*kernel[7]+tmp[4675]*kernel[8];
				ans[4575]<=tmp[4474]*kernel[0]+tmp[4475]*kernel[1]+tmp[4476]*kernel[2]+tmp[4574]*kernel[3]+tmp[4575]*kernel[4]+tmp[4576]*kernel[5]+tmp[4674]*kernel[6]+tmp[4675]*kernel[7]+tmp[4676]*kernel[8];
				ans[4576]<=tmp[4475]*kernel[0]+tmp[4476]*kernel[1]+tmp[4477]*kernel[2]+tmp[4575]*kernel[3]+tmp[4576]*kernel[4]+tmp[4577]*kernel[5]+tmp[4675]*kernel[6]+tmp[4676]*kernel[7]+tmp[4677]*kernel[8];
				ans[4577]<=tmp[4476]*kernel[0]+tmp[4477]*kernel[1]+tmp[4478]*kernel[2]+tmp[4576]*kernel[3]+tmp[4577]*kernel[4]+tmp[4578]*kernel[5]+tmp[4676]*kernel[6]+tmp[4677]*kernel[7]+tmp[4678]*kernel[8];
				ans[4578]<=tmp[4477]*kernel[0]+tmp[4478]*kernel[1]+tmp[4479]*kernel[2]+tmp[4577]*kernel[3]+tmp[4578]*kernel[4]+tmp[4579]*kernel[5]+tmp[4677]*kernel[6]+tmp[4678]*kernel[7]+tmp[4679]*kernel[8];
				ans[4579]<=tmp[4478]*kernel[0]+tmp[4479]*kernel[1]+tmp[4480]*kernel[2]+tmp[4578]*kernel[3]+tmp[4579]*kernel[4]+tmp[4580]*kernel[5]+tmp[4678]*kernel[6]+tmp[4679]*kernel[7]+tmp[4680]*kernel[8];
				ans[4580]<=tmp[4479]*kernel[0]+tmp[4480]*kernel[1]+tmp[4481]*kernel[2]+tmp[4579]*kernel[3]+tmp[4580]*kernel[4]+tmp[4581]*kernel[5]+tmp[4679]*kernel[6]+tmp[4680]*kernel[7]+tmp[4681]*kernel[8];
				ans[4581]<=tmp[4480]*kernel[0]+tmp[4481]*kernel[1]+tmp[4482]*kernel[2]+tmp[4580]*kernel[3]+tmp[4581]*kernel[4]+tmp[4582]*kernel[5]+tmp[4680]*kernel[6]+tmp[4681]*kernel[7]+tmp[4682]*kernel[8];
				ans[4582]<=tmp[4481]*kernel[0]+tmp[4482]*kernel[1]+tmp[4483]*kernel[2]+tmp[4581]*kernel[3]+tmp[4582]*kernel[4]+tmp[4583]*kernel[5]+tmp[4681]*kernel[6]+tmp[4682]*kernel[7]+tmp[4683]*kernel[8];
				ans[4583]<=tmp[4482]*kernel[0]+tmp[4483]*kernel[1]+tmp[4484]*kernel[2]+tmp[4582]*kernel[3]+tmp[4583]*kernel[4]+tmp[4584]*kernel[5]+tmp[4682]*kernel[6]+tmp[4683]*kernel[7]+tmp[4684]*kernel[8];
				ans[4584]<=tmp[4483]*kernel[0]+tmp[4484]*kernel[1]+tmp[4485]*kernel[2]+tmp[4583]*kernel[3]+tmp[4584]*kernel[4]+tmp[4585]*kernel[5]+tmp[4683]*kernel[6]+tmp[4684]*kernel[7]+tmp[4685]*kernel[8];
				ans[4585]<=tmp[4484]*kernel[0]+tmp[4485]*kernel[1]+tmp[4486]*kernel[2]+tmp[4584]*kernel[3]+tmp[4585]*kernel[4]+tmp[4586]*kernel[5]+tmp[4684]*kernel[6]+tmp[4685]*kernel[7]+tmp[4686]*kernel[8];
				ans[4586]<=tmp[4485]*kernel[0]+tmp[4486]*kernel[1]+tmp[4487]*kernel[2]+tmp[4585]*kernel[3]+tmp[4586]*kernel[4]+tmp[4587]*kernel[5]+tmp[4685]*kernel[6]+tmp[4686]*kernel[7]+tmp[4687]*kernel[8];
				ans[4587]<=tmp[4486]*kernel[0]+tmp[4487]*kernel[1]+tmp[4488]*kernel[2]+tmp[4586]*kernel[3]+tmp[4587]*kernel[4]+tmp[4588]*kernel[5]+tmp[4686]*kernel[6]+tmp[4687]*kernel[7]+tmp[4688]*kernel[8];
				ans[4588]<=tmp[4487]*kernel[0]+tmp[4488]*kernel[1]+tmp[4489]*kernel[2]+tmp[4587]*kernel[3]+tmp[4588]*kernel[4]+tmp[4589]*kernel[5]+tmp[4687]*kernel[6]+tmp[4688]*kernel[7]+tmp[4689]*kernel[8];
				ans[4589]<=tmp[4488]*kernel[0]+tmp[4489]*kernel[1]+tmp[4490]*kernel[2]+tmp[4588]*kernel[3]+tmp[4589]*kernel[4]+tmp[4590]*kernel[5]+tmp[4688]*kernel[6]+tmp[4689]*kernel[7]+tmp[4690]*kernel[8];
				ans[4590]<=tmp[4489]*kernel[0]+tmp[4490]*kernel[1]+tmp[4491]*kernel[2]+tmp[4589]*kernel[3]+tmp[4590]*kernel[4]+tmp[4591]*kernel[5]+tmp[4689]*kernel[6]+tmp[4690]*kernel[7]+tmp[4691]*kernel[8];
				ans[4591]<=tmp[4490]*kernel[0]+tmp[4491]*kernel[1]+tmp[4492]*kernel[2]+tmp[4590]*kernel[3]+tmp[4591]*kernel[4]+tmp[4592]*kernel[5]+tmp[4690]*kernel[6]+tmp[4691]*kernel[7]+tmp[4692]*kernel[8];
				ans[4592]<=tmp[4491]*kernel[0]+tmp[4492]*kernel[1]+tmp[4493]*kernel[2]+tmp[4591]*kernel[3]+tmp[4592]*kernel[4]+tmp[4593]*kernel[5]+tmp[4691]*kernel[6]+tmp[4692]*kernel[7]+tmp[4693]*kernel[8];
				ans[4593]<=tmp[4492]*kernel[0]+tmp[4493]*kernel[1]+tmp[4494]*kernel[2]+tmp[4592]*kernel[3]+tmp[4593]*kernel[4]+tmp[4594]*kernel[5]+tmp[4692]*kernel[6]+tmp[4693]*kernel[7]+tmp[4694]*kernel[8];
				ans[4594]<=tmp[4493]*kernel[0]+tmp[4494]*kernel[1]+tmp[4495]*kernel[2]+tmp[4593]*kernel[3]+tmp[4594]*kernel[4]+tmp[4595]*kernel[5]+tmp[4693]*kernel[6]+tmp[4694]*kernel[7]+tmp[4695]*kernel[8];
				ans[4595]<=tmp[4494]*kernel[0]+tmp[4495]*kernel[1]+tmp[4496]*kernel[2]+tmp[4594]*kernel[3]+tmp[4595]*kernel[4]+tmp[4596]*kernel[5]+tmp[4694]*kernel[6]+tmp[4695]*kernel[7]+tmp[4696]*kernel[8];
				ans[4596]<=tmp[4495]*kernel[0]+tmp[4496]*kernel[1]+tmp[4497]*kernel[2]+tmp[4595]*kernel[3]+tmp[4596]*kernel[4]+tmp[4597]*kernel[5]+tmp[4695]*kernel[6]+tmp[4696]*kernel[7]+tmp[4697]*kernel[8];
				ans[4597]<=tmp[4496]*kernel[0]+tmp[4497]*kernel[1]+tmp[4498]*kernel[2]+tmp[4596]*kernel[3]+tmp[4597]*kernel[4]+tmp[4598]*kernel[5]+tmp[4696]*kernel[6]+tmp[4697]*kernel[7]+tmp[4698]*kernel[8];
				ans[4598]<=tmp[4497]*kernel[0]+tmp[4498]*kernel[1]+tmp[4499]*kernel[2]+tmp[4597]*kernel[3]+tmp[4598]*kernel[4]+tmp[4599]*kernel[5]+tmp[4697]*kernel[6]+tmp[4698]*kernel[7]+tmp[4699]*kernel[8];
				ans[4599]<=tmp[4498]*kernel[0]+tmp[4499]*kernel[1]+tmp[4598]*kernel[3]+tmp[4599]*kernel[4]+tmp[4698]*kernel[6]+tmp[4699]*kernel[7];
				ans[4600]<=tmp[4500]*kernel[1]+tmp[4501]*kernel[2]+tmp[4600]*kernel[4]+tmp[4601]*kernel[5]+tmp[4700]*kernel[7]+tmp[4701]*kernel[8];
				ans[4601]<=tmp[4500]*kernel[0]+tmp[4501]*kernel[1]+tmp[4502]*kernel[2]+tmp[4600]*kernel[3]+tmp[4601]*kernel[4]+tmp[4602]*kernel[5]+tmp[4700]*kernel[6]+tmp[4701]*kernel[7]+tmp[4702]*kernel[8];
				ans[4602]<=tmp[4501]*kernel[0]+tmp[4502]*kernel[1]+tmp[4503]*kernel[2]+tmp[4601]*kernel[3]+tmp[4602]*kernel[4]+tmp[4603]*kernel[5]+tmp[4701]*kernel[6]+tmp[4702]*kernel[7]+tmp[4703]*kernel[8];
				ans[4603]<=tmp[4502]*kernel[0]+tmp[4503]*kernel[1]+tmp[4504]*kernel[2]+tmp[4602]*kernel[3]+tmp[4603]*kernel[4]+tmp[4604]*kernel[5]+tmp[4702]*kernel[6]+tmp[4703]*kernel[7]+tmp[4704]*kernel[8];
				ans[4604]<=tmp[4503]*kernel[0]+tmp[4504]*kernel[1]+tmp[4505]*kernel[2]+tmp[4603]*kernel[3]+tmp[4604]*kernel[4]+tmp[4605]*kernel[5]+tmp[4703]*kernel[6]+tmp[4704]*kernel[7]+tmp[4705]*kernel[8];
				ans[4605]<=tmp[4504]*kernel[0]+tmp[4505]*kernel[1]+tmp[4506]*kernel[2]+tmp[4604]*kernel[3]+tmp[4605]*kernel[4]+tmp[4606]*kernel[5]+tmp[4704]*kernel[6]+tmp[4705]*kernel[7]+tmp[4706]*kernel[8];
				ans[4606]<=tmp[4505]*kernel[0]+tmp[4506]*kernel[1]+tmp[4507]*kernel[2]+tmp[4605]*kernel[3]+tmp[4606]*kernel[4]+tmp[4607]*kernel[5]+tmp[4705]*kernel[6]+tmp[4706]*kernel[7]+tmp[4707]*kernel[8];
				ans[4607]<=tmp[4506]*kernel[0]+tmp[4507]*kernel[1]+tmp[4508]*kernel[2]+tmp[4606]*kernel[3]+tmp[4607]*kernel[4]+tmp[4608]*kernel[5]+tmp[4706]*kernel[6]+tmp[4707]*kernel[7]+tmp[4708]*kernel[8];
				ans[4608]<=tmp[4507]*kernel[0]+tmp[4508]*kernel[1]+tmp[4509]*kernel[2]+tmp[4607]*kernel[3]+tmp[4608]*kernel[4]+tmp[4609]*kernel[5]+tmp[4707]*kernel[6]+tmp[4708]*kernel[7]+tmp[4709]*kernel[8];
				ans[4609]<=tmp[4508]*kernel[0]+tmp[4509]*kernel[1]+tmp[4510]*kernel[2]+tmp[4608]*kernel[3]+tmp[4609]*kernel[4]+tmp[4610]*kernel[5]+tmp[4708]*kernel[6]+tmp[4709]*kernel[7]+tmp[4710]*kernel[8];
				ans[4610]<=tmp[4509]*kernel[0]+tmp[4510]*kernel[1]+tmp[4511]*kernel[2]+tmp[4609]*kernel[3]+tmp[4610]*kernel[4]+tmp[4611]*kernel[5]+tmp[4709]*kernel[6]+tmp[4710]*kernel[7]+tmp[4711]*kernel[8];
				ans[4611]<=tmp[4510]*kernel[0]+tmp[4511]*kernel[1]+tmp[4512]*kernel[2]+tmp[4610]*kernel[3]+tmp[4611]*kernel[4]+tmp[4612]*kernel[5]+tmp[4710]*kernel[6]+tmp[4711]*kernel[7]+tmp[4712]*kernel[8];
				ans[4612]<=tmp[4511]*kernel[0]+tmp[4512]*kernel[1]+tmp[4513]*kernel[2]+tmp[4611]*kernel[3]+tmp[4612]*kernel[4]+tmp[4613]*kernel[5]+tmp[4711]*kernel[6]+tmp[4712]*kernel[7]+tmp[4713]*kernel[8];
				ans[4613]<=tmp[4512]*kernel[0]+tmp[4513]*kernel[1]+tmp[4514]*kernel[2]+tmp[4612]*kernel[3]+tmp[4613]*kernel[4]+tmp[4614]*kernel[5]+tmp[4712]*kernel[6]+tmp[4713]*kernel[7]+tmp[4714]*kernel[8];
				ans[4614]<=tmp[4513]*kernel[0]+tmp[4514]*kernel[1]+tmp[4515]*kernel[2]+tmp[4613]*kernel[3]+tmp[4614]*kernel[4]+tmp[4615]*kernel[5]+tmp[4713]*kernel[6]+tmp[4714]*kernel[7]+tmp[4715]*kernel[8];
				ans[4615]<=tmp[4514]*kernel[0]+tmp[4515]*kernel[1]+tmp[4516]*kernel[2]+tmp[4614]*kernel[3]+tmp[4615]*kernel[4]+tmp[4616]*kernel[5]+tmp[4714]*kernel[6]+tmp[4715]*kernel[7]+tmp[4716]*kernel[8];
				ans[4616]<=tmp[4515]*kernel[0]+tmp[4516]*kernel[1]+tmp[4517]*kernel[2]+tmp[4615]*kernel[3]+tmp[4616]*kernel[4]+tmp[4617]*kernel[5]+tmp[4715]*kernel[6]+tmp[4716]*kernel[7]+tmp[4717]*kernel[8];
				ans[4617]<=tmp[4516]*kernel[0]+tmp[4517]*kernel[1]+tmp[4518]*kernel[2]+tmp[4616]*kernel[3]+tmp[4617]*kernel[4]+tmp[4618]*kernel[5]+tmp[4716]*kernel[6]+tmp[4717]*kernel[7]+tmp[4718]*kernel[8];
				ans[4618]<=tmp[4517]*kernel[0]+tmp[4518]*kernel[1]+tmp[4519]*kernel[2]+tmp[4617]*kernel[3]+tmp[4618]*kernel[4]+tmp[4619]*kernel[5]+tmp[4717]*kernel[6]+tmp[4718]*kernel[7]+tmp[4719]*kernel[8];
				ans[4619]<=tmp[4518]*kernel[0]+tmp[4519]*kernel[1]+tmp[4520]*kernel[2]+tmp[4618]*kernel[3]+tmp[4619]*kernel[4]+tmp[4620]*kernel[5]+tmp[4718]*kernel[6]+tmp[4719]*kernel[7]+tmp[4720]*kernel[8];
				ans[4620]<=tmp[4519]*kernel[0]+tmp[4520]*kernel[1]+tmp[4521]*kernel[2]+tmp[4619]*kernel[3]+tmp[4620]*kernel[4]+tmp[4621]*kernel[5]+tmp[4719]*kernel[6]+tmp[4720]*kernel[7]+tmp[4721]*kernel[8];
				ans[4621]<=tmp[4520]*kernel[0]+tmp[4521]*kernel[1]+tmp[4522]*kernel[2]+tmp[4620]*kernel[3]+tmp[4621]*kernel[4]+tmp[4622]*kernel[5]+tmp[4720]*kernel[6]+tmp[4721]*kernel[7]+tmp[4722]*kernel[8];
				ans[4622]<=tmp[4521]*kernel[0]+tmp[4522]*kernel[1]+tmp[4523]*kernel[2]+tmp[4621]*kernel[3]+tmp[4622]*kernel[4]+tmp[4623]*kernel[5]+tmp[4721]*kernel[6]+tmp[4722]*kernel[7]+tmp[4723]*kernel[8];
				ans[4623]<=tmp[4522]*kernel[0]+tmp[4523]*kernel[1]+tmp[4524]*kernel[2]+tmp[4622]*kernel[3]+tmp[4623]*kernel[4]+tmp[4624]*kernel[5]+tmp[4722]*kernel[6]+tmp[4723]*kernel[7]+tmp[4724]*kernel[8];
				ans[4624]<=tmp[4523]*kernel[0]+tmp[4524]*kernel[1]+tmp[4525]*kernel[2]+tmp[4623]*kernel[3]+tmp[4624]*kernel[4]+tmp[4625]*kernel[5]+tmp[4723]*kernel[6]+tmp[4724]*kernel[7]+tmp[4725]*kernel[8];
				ans[4625]<=tmp[4524]*kernel[0]+tmp[4525]*kernel[1]+tmp[4526]*kernel[2]+tmp[4624]*kernel[3]+tmp[4625]*kernel[4]+tmp[4626]*kernel[5]+tmp[4724]*kernel[6]+tmp[4725]*kernel[7]+tmp[4726]*kernel[8];
				ans[4626]<=tmp[4525]*kernel[0]+tmp[4526]*kernel[1]+tmp[4527]*kernel[2]+tmp[4625]*kernel[3]+tmp[4626]*kernel[4]+tmp[4627]*kernel[5]+tmp[4725]*kernel[6]+tmp[4726]*kernel[7]+tmp[4727]*kernel[8];
				ans[4627]<=tmp[4526]*kernel[0]+tmp[4527]*kernel[1]+tmp[4528]*kernel[2]+tmp[4626]*kernel[3]+tmp[4627]*kernel[4]+tmp[4628]*kernel[5]+tmp[4726]*kernel[6]+tmp[4727]*kernel[7]+tmp[4728]*kernel[8];
				ans[4628]<=tmp[4527]*kernel[0]+tmp[4528]*kernel[1]+tmp[4529]*kernel[2]+tmp[4627]*kernel[3]+tmp[4628]*kernel[4]+tmp[4629]*kernel[5]+tmp[4727]*kernel[6]+tmp[4728]*kernel[7]+tmp[4729]*kernel[8];
				ans[4629]<=tmp[4528]*kernel[0]+tmp[4529]*kernel[1]+tmp[4530]*kernel[2]+tmp[4628]*kernel[3]+tmp[4629]*kernel[4]+tmp[4630]*kernel[5]+tmp[4728]*kernel[6]+tmp[4729]*kernel[7]+tmp[4730]*kernel[8];
				ans[4630]<=tmp[4529]*kernel[0]+tmp[4530]*kernel[1]+tmp[4531]*kernel[2]+tmp[4629]*kernel[3]+tmp[4630]*kernel[4]+tmp[4631]*kernel[5]+tmp[4729]*kernel[6]+tmp[4730]*kernel[7]+tmp[4731]*kernel[8];
				ans[4631]<=tmp[4530]*kernel[0]+tmp[4531]*kernel[1]+tmp[4532]*kernel[2]+tmp[4630]*kernel[3]+tmp[4631]*kernel[4]+tmp[4632]*kernel[5]+tmp[4730]*kernel[6]+tmp[4731]*kernel[7]+tmp[4732]*kernel[8];
				ans[4632]<=tmp[4531]*kernel[0]+tmp[4532]*kernel[1]+tmp[4533]*kernel[2]+tmp[4631]*kernel[3]+tmp[4632]*kernel[4]+tmp[4633]*kernel[5]+tmp[4731]*kernel[6]+tmp[4732]*kernel[7]+tmp[4733]*kernel[8];
				ans[4633]<=tmp[4532]*kernel[0]+tmp[4533]*kernel[1]+tmp[4534]*kernel[2]+tmp[4632]*kernel[3]+tmp[4633]*kernel[4]+tmp[4634]*kernel[5]+tmp[4732]*kernel[6]+tmp[4733]*kernel[7]+tmp[4734]*kernel[8];
				ans[4634]<=tmp[4533]*kernel[0]+tmp[4534]*kernel[1]+tmp[4535]*kernel[2]+tmp[4633]*kernel[3]+tmp[4634]*kernel[4]+tmp[4635]*kernel[5]+tmp[4733]*kernel[6]+tmp[4734]*kernel[7]+tmp[4735]*kernel[8];
				ans[4635]<=tmp[4534]*kernel[0]+tmp[4535]*kernel[1]+tmp[4536]*kernel[2]+tmp[4634]*kernel[3]+tmp[4635]*kernel[4]+tmp[4636]*kernel[5]+tmp[4734]*kernel[6]+tmp[4735]*kernel[7]+tmp[4736]*kernel[8];
				ans[4636]<=tmp[4535]*kernel[0]+tmp[4536]*kernel[1]+tmp[4537]*kernel[2]+tmp[4635]*kernel[3]+tmp[4636]*kernel[4]+tmp[4637]*kernel[5]+tmp[4735]*kernel[6]+tmp[4736]*kernel[7]+tmp[4737]*kernel[8];
				ans[4637]<=tmp[4536]*kernel[0]+tmp[4537]*kernel[1]+tmp[4538]*kernel[2]+tmp[4636]*kernel[3]+tmp[4637]*kernel[4]+tmp[4638]*kernel[5]+tmp[4736]*kernel[6]+tmp[4737]*kernel[7]+tmp[4738]*kernel[8];
				ans[4638]<=tmp[4537]*kernel[0]+tmp[4538]*kernel[1]+tmp[4539]*kernel[2]+tmp[4637]*kernel[3]+tmp[4638]*kernel[4]+tmp[4639]*kernel[5]+tmp[4737]*kernel[6]+tmp[4738]*kernel[7]+tmp[4739]*kernel[8];
				ans[4639]<=tmp[4538]*kernel[0]+tmp[4539]*kernel[1]+tmp[4540]*kernel[2]+tmp[4638]*kernel[3]+tmp[4639]*kernel[4]+tmp[4640]*kernel[5]+tmp[4738]*kernel[6]+tmp[4739]*kernel[7]+tmp[4740]*kernel[8];
				ans[4640]<=tmp[4539]*kernel[0]+tmp[4540]*kernel[1]+tmp[4541]*kernel[2]+tmp[4639]*kernel[3]+tmp[4640]*kernel[4]+tmp[4641]*kernel[5]+tmp[4739]*kernel[6]+tmp[4740]*kernel[7]+tmp[4741]*kernel[8];
				ans[4641]<=tmp[4540]*kernel[0]+tmp[4541]*kernel[1]+tmp[4542]*kernel[2]+tmp[4640]*kernel[3]+tmp[4641]*kernel[4]+tmp[4642]*kernel[5]+tmp[4740]*kernel[6]+tmp[4741]*kernel[7]+tmp[4742]*kernel[8];
				ans[4642]<=tmp[4541]*kernel[0]+tmp[4542]*kernel[1]+tmp[4543]*kernel[2]+tmp[4641]*kernel[3]+tmp[4642]*kernel[4]+tmp[4643]*kernel[5]+tmp[4741]*kernel[6]+tmp[4742]*kernel[7]+tmp[4743]*kernel[8];
				ans[4643]<=tmp[4542]*kernel[0]+tmp[4543]*kernel[1]+tmp[4544]*kernel[2]+tmp[4642]*kernel[3]+tmp[4643]*kernel[4]+tmp[4644]*kernel[5]+tmp[4742]*kernel[6]+tmp[4743]*kernel[7]+tmp[4744]*kernel[8];
				ans[4644]<=tmp[4543]*kernel[0]+tmp[4544]*kernel[1]+tmp[4545]*kernel[2]+tmp[4643]*kernel[3]+tmp[4644]*kernel[4]+tmp[4645]*kernel[5]+tmp[4743]*kernel[6]+tmp[4744]*kernel[7]+tmp[4745]*kernel[8];
				ans[4645]<=tmp[4544]*kernel[0]+tmp[4545]*kernel[1]+tmp[4546]*kernel[2]+tmp[4644]*kernel[3]+tmp[4645]*kernel[4]+tmp[4646]*kernel[5]+tmp[4744]*kernel[6]+tmp[4745]*kernel[7]+tmp[4746]*kernel[8];
				ans[4646]<=tmp[4545]*kernel[0]+tmp[4546]*kernel[1]+tmp[4547]*kernel[2]+tmp[4645]*kernel[3]+tmp[4646]*kernel[4]+tmp[4647]*kernel[5]+tmp[4745]*kernel[6]+tmp[4746]*kernel[7]+tmp[4747]*kernel[8];
				ans[4647]<=tmp[4546]*kernel[0]+tmp[4547]*kernel[1]+tmp[4548]*kernel[2]+tmp[4646]*kernel[3]+tmp[4647]*kernel[4]+tmp[4648]*kernel[5]+tmp[4746]*kernel[6]+tmp[4747]*kernel[7]+tmp[4748]*kernel[8];
				ans[4648]<=tmp[4547]*kernel[0]+tmp[4548]*kernel[1]+tmp[4549]*kernel[2]+tmp[4647]*kernel[3]+tmp[4648]*kernel[4]+tmp[4649]*kernel[5]+tmp[4747]*kernel[6]+tmp[4748]*kernel[7]+tmp[4749]*kernel[8];
				ans[4649]<=tmp[4548]*kernel[0]+tmp[4549]*kernel[1]+tmp[4550]*kernel[2]+tmp[4648]*kernel[3]+tmp[4649]*kernel[4]+tmp[4650]*kernel[5]+tmp[4748]*kernel[6]+tmp[4749]*kernel[7]+tmp[4750]*kernel[8];
				ans[4650]<=tmp[4549]*kernel[0]+tmp[4550]*kernel[1]+tmp[4551]*kernel[2]+tmp[4649]*kernel[3]+tmp[4650]*kernel[4]+tmp[4651]*kernel[5]+tmp[4749]*kernel[6]+tmp[4750]*kernel[7]+tmp[4751]*kernel[8];
				ans[4651]<=tmp[4550]*kernel[0]+tmp[4551]*kernel[1]+tmp[4552]*kernel[2]+tmp[4650]*kernel[3]+tmp[4651]*kernel[4]+tmp[4652]*kernel[5]+tmp[4750]*kernel[6]+tmp[4751]*kernel[7]+tmp[4752]*kernel[8];
				ans[4652]<=tmp[4551]*kernel[0]+tmp[4552]*kernel[1]+tmp[4553]*kernel[2]+tmp[4651]*kernel[3]+tmp[4652]*kernel[4]+tmp[4653]*kernel[5]+tmp[4751]*kernel[6]+tmp[4752]*kernel[7]+tmp[4753]*kernel[8];
				ans[4653]<=tmp[4552]*kernel[0]+tmp[4553]*kernel[1]+tmp[4554]*kernel[2]+tmp[4652]*kernel[3]+tmp[4653]*kernel[4]+tmp[4654]*kernel[5]+tmp[4752]*kernel[6]+tmp[4753]*kernel[7]+tmp[4754]*kernel[8];
				ans[4654]<=tmp[4553]*kernel[0]+tmp[4554]*kernel[1]+tmp[4555]*kernel[2]+tmp[4653]*kernel[3]+tmp[4654]*kernel[4]+tmp[4655]*kernel[5]+tmp[4753]*kernel[6]+tmp[4754]*kernel[7]+tmp[4755]*kernel[8];
				ans[4655]<=tmp[4554]*kernel[0]+tmp[4555]*kernel[1]+tmp[4556]*kernel[2]+tmp[4654]*kernel[3]+tmp[4655]*kernel[4]+tmp[4656]*kernel[5]+tmp[4754]*kernel[6]+tmp[4755]*kernel[7]+tmp[4756]*kernel[8];
				ans[4656]<=tmp[4555]*kernel[0]+tmp[4556]*kernel[1]+tmp[4557]*kernel[2]+tmp[4655]*kernel[3]+tmp[4656]*kernel[4]+tmp[4657]*kernel[5]+tmp[4755]*kernel[6]+tmp[4756]*kernel[7]+tmp[4757]*kernel[8];
				ans[4657]<=tmp[4556]*kernel[0]+tmp[4557]*kernel[1]+tmp[4558]*kernel[2]+tmp[4656]*kernel[3]+tmp[4657]*kernel[4]+tmp[4658]*kernel[5]+tmp[4756]*kernel[6]+tmp[4757]*kernel[7]+tmp[4758]*kernel[8];
				ans[4658]<=tmp[4557]*kernel[0]+tmp[4558]*kernel[1]+tmp[4559]*kernel[2]+tmp[4657]*kernel[3]+tmp[4658]*kernel[4]+tmp[4659]*kernel[5]+tmp[4757]*kernel[6]+tmp[4758]*kernel[7]+tmp[4759]*kernel[8];
				ans[4659]<=tmp[4558]*kernel[0]+tmp[4559]*kernel[1]+tmp[4560]*kernel[2]+tmp[4658]*kernel[3]+tmp[4659]*kernel[4]+tmp[4660]*kernel[5]+tmp[4758]*kernel[6]+tmp[4759]*kernel[7]+tmp[4760]*kernel[8];
				ans[4660]<=tmp[4559]*kernel[0]+tmp[4560]*kernel[1]+tmp[4561]*kernel[2]+tmp[4659]*kernel[3]+tmp[4660]*kernel[4]+tmp[4661]*kernel[5]+tmp[4759]*kernel[6]+tmp[4760]*kernel[7]+tmp[4761]*kernel[8];
				ans[4661]<=tmp[4560]*kernel[0]+tmp[4561]*kernel[1]+tmp[4562]*kernel[2]+tmp[4660]*kernel[3]+tmp[4661]*kernel[4]+tmp[4662]*kernel[5]+tmp[4760]*kernel[6]+tmp[4761]*kernel[7]+tmp[4762]*kernel[8];
				ans[4662]<=tmp[4561]*kernel[0]+tmp[4562]*kernel[1]+tmp[4563]*kernel[2]+tmp[4661]*kernel[3]+tmp[4662]*kernel[4]+tmp[4663]*kernel[5]+tmp[4761]*kernel[6]+tmp[4762]*kernel[7]+tmp[4763]*kernel[8];
				ans[4663]<=tmp[4562]*kernel[0]+tmp[4563]*kernel[1]+tmp[4564]*kernel[2]+tmp[4662]*kernel[3]+tmp[4663]*kernel[4]+tmp[4664]*kernel[5]+tmp[4762]*kernel[6]+tmp[4763]*kernel[7]+tmp[4764]*kernel[8];
				ans[4664]<=tmp[4563]*kernel[0]+tmp[4564]*kernel[1]+tmp[4565]*kernel[2]+tmp[4663]*kernel[3]+tmp[4664]*kernel[4]+tmp[4665]*kernel[5]+tmp[4763]*kernel[6]+tmp[4764]*kernel[7]+tmp[4765]*kernel[8];
				ans[4665]<=tmp[4564]*kernel[0]+tmp[4565]*kernel[1]+tmp[4566]*kernel[2]+tmp[4664]*kernel[3]+tmp[4665]*kernel[4]+tmp[4666]*kernel[5]+tmp[4764]*kernel[6]+tmp[4765]*kernel[7]+tmp[4766]*kernel[8];
				ans[4666]<=tmp[4565]*kernel[0]+tmp[4566]*kernel[1]+tmp[4567]*kernel[2]+tmp[4665]*kernel[3]+tmp[4666]*kernel[4]+tmp[4667]*kernel[5]+tmp[4765]*kernel[6]+tmp[4766]*kernel[7]+tmp[4767]*kernel[8];
				ans[4667]<=tmp[4566]*kernel[0]+tmp[4567]*kernel[1]+tmp[4568]*kernel[2]+tmp[4666]*kernel[3]+tmp[4667]*kernel[4]+tmp[4668]*kernel[5]+tmp[4766]*kernel[6]+tmp[4767]*kernel[7]+tmp[4768]*kernel[8];
				ans[4668]<=tmp[4567]*kernel[0]+tmp[4568]*kernel[1]+tmp[4569]*kernel[2]+tmp[4667]*kernel[3]+tmp[4668]*kernel[4]+tmp[4669]*kernel[5]+tmp[4767]*kernel[6]+tmp[4768]*kernel[7]+tmp[4769]*kernel[8];
				ans[4669]<=tmp[4568]*kernel[0]+tmp[4569]*kernel[1]+tmp[4570]*kernel[2]+tmp[4668]*kernel[3]+tmp[4669]*kernel[4]+tmp[4670]*kernel[5]+tmp[4768]*kernel[6]+tmp[4769]*kernel[7]+tmp[4770]*kernel[8];
				ans[4670]<=tmp[4569]*kernel[0]+tmp[4570]*kernel[1]+tmp[4571]*kernel[2]+tmp[4669]*kernel[3]+tmp[4670]*kernel[4]+tmp[4671]*kernel[5]+tmp[4769]*kernel[6]+tmp[4770]*kernel[7]+tmp[4771]*kernel[8];
				ans[4671]<=tmp[4570]*kernel[0]+tmp[4571]*kernel[1]+tmp[4572]*kernel[2]+tmp[4670]*kernel[3]+tmp[4671]*kernel[4]+tmp[4672]*kernel[5]+tmp[4770]*kernel[6]+tmp[4771]*kernel[7]+tmp[4772]*kernel[8];
				ans[4672]<=tmp[4571]*kernel[0]+tmp[4572]*kernel[1]+tmp[4573]*kernel[2]+tmp[4671]*kernel[3]+tmp[4672]*kernel[4]+tmp[4673]*kernel[5]+tmp[4771]*kernel[6]+tmp[4772]*kernel[7]+tmp[4773]*kernel[8];
				ans[4673]<=tmp[4572]*kernel[0]+tmp[4573]*kernel[1]+tmp[4574]*kernel[2]+tmp[4672]*kernel[3]+tmp[4673]*kernel[4]+tmp[4674]*kernel[5]+tmp[4772]*kernel[6]+tmp[4773]*kernel[7]+tmp[4774]*kernel[8];
				ans[4674]<=tmp[4573]*kernel[0]+tmp[4574]*kernel[1]+tmp[4575]*kernel[2]+tmp[4673]*kernel[3]+tmp[4674]*kernel[4]+tmp[4675]*kernel[5]+tmp[4773]*kernel[6]+tmp[4774]*kernel[7]+tmp[4775]*kernel[8];
				ans[4675]<=tmp[4574]*kernel[0]+tmp[4575]*kernel[1]+tmp[4576]*kernel[2]+tmp[4674]*kernel[3]+tmp[4675]*kernel[4]+tmp[4676]*kernel[5]+tmp[4774]*kernel[6]+tmp[4775]*kernel[7]+tmp[4776]*kernel[8];
				ans[4676]<=tmp[4575]*kernel[0]+tmp[4576]*kernel[1]+tmp[4577]*kernel[2]+tmp[4675]*kernel[3]+tmp[4676]*kernel[4]+tmp[4677]*kernel[5]+tmp[4775]*kernel[6]+tmp[4776]*kernel[7]+tmp[4777]*kernel[8];
				ans[4677]<=tmp[4576]*kernel[0]+tmp[4577]*kernel[1]+tmp[4578]*kernel[2]+tmp[4676]*kernel[3]+tmp[4677]*kernel[4]+tmp[4678]*kernel[5]+tmp[4776]*kernel[6]+tmp[4777]*kernel[7]+tmp[4778]*kernel[8];
				ans[4678]<=tmp[4577]*kernel[0]+tmp[4578]*kernel[1]+tmp[4579]*kernel[2]+tmp[4677]*kernel[3]+tmp[4678]*kernel[4]+tmp[4679]*kernel[5]+tmp[4777]*kernel[6]+tmp[4778]*kernel[7]+tmp[4779]*kernel[8];
				ans[4679]<=tmp[4578]*kernel[0]+tmp[4579]*kernel[1]+tmp[4580]*kernel[2]+tmp[4678]*kernel[3]+tmp[4679]*kernel[4]+tmp[4680]*kernel[5]+tmp[4778]*kernel[6]+tmp[4779]*kernel[7]+tmp[4780]*kernel[8];
				ans[4680]<=tmp[4579]*kernel[0]+tmp[4580]*kernel[1]+tmp[4581]*kernel[2]+tmp[4679]*kernel[3]+tmp[4680]*kernel[4]+tmp[4681]*kernel[5]+tmp[4779]*kernel[6]+tmp[4780]*kernel[7]+tmp[4781]*kernel[8];
				ans[4681]<=tmp[4580]*kernel[0]+tmp[4581]*kernel[1]+tmp[4582]*kernel[2]+tmp[4680]*kernel[3]+tmp[4681]*kernel[4]+tmp[4682]*kernel[5]+tmp[4780]*kernel[6]+tmp[4781]*kernel[7]+tmp[4782]*kernel[8];
				ans[4682]<=tmp[4581]*kernel[0]+tmp[4582]*kernel[1]+tmp[4583]*kernel[2]+tmp[4681]*kernel[3]+tmp[4682]*kernel[4]+tmp[4683]*kernel[5]+tmp[4781]*kernel[6]+tmp[4782]*kernel[7]+tmp[4783]*kernel[8];
				ans[4683]<=tmp[4582]*kernel[0]+tmp[4583]*kernel[1]+tmp[4584]*kernel[2]+tmp[4682]*kernel[3]+tmp[4683]*kernel[4]+tmp[4684]*kernel[5]+tmp[4782]*kernel[6]+tmp[4783]*kernel[7]+tmp[4784]*kernel[8];
				ans[4684]<=tmp[4583]*kernel[0]+tmp[4584]*kernel[1]+tmp[4585]*kernel[2]+tmp[4683]*kernel[3]+tmp[4684]*kernel[4]+tmp[4685]*kernel[5]+tmp[4783]*kernel[6]+tmp[4784]*kernel[7]+tmp[4785]*kernel[8];
				ans[4685]<=tmp[4584]*kernel[0]+tmp[4585]*kernel[1]+tmp[4586]*kernel[2]+tmp[4684]*kernel[3]+tmp[4685]*kernel[4]+tmp[4686]*kernel[5]+tmp[4784]*kernel[6]+tmp[4785]*kernel[7]+tmp[4786]*kernel[8];
				ans[4686]<=tmp[4585]*kernel[0]+tmp[4586]*kernel[1]+tmp[4587]*kernel[2]+tmp[4685]*kernel[3]+tmp[4686]*kernel[4]+tmp[4687]*kernel[5]+tmp[4785]*kernel[6]+tmp[4786]*kernel[7]+tmp[4787]*kernel[8];
				ans[4687]<=tmp[4586]*kernel[0]+tmp[4587]*kernel[1]+tmp[4588]*kernel[2]+tmp[4686]*kernel[3]+tmp[4687]*kernel[4]+tmp[4688]*kernel[5]+tmp[4786]*kernel[6]+tmp[4787]*kernel[7]+tmp[4788]*kernel[8];
				ans[4688]<=tmp[4587]*kernel[0]+tmp[4588]*kernel[1]+tmp[4589]*kernel[2]+tmp[4687]*kernel[3]+tmp[4688]*kernel[4]+tmp[4689]*kernel[5]+tmp[4787]*kernel[6]+tmp[4788]*kernel[7]+tmp[4789]*kernel[8];
				ans[4689]<=tmp[4588]*kernel[0]+tmp[4589]*kernel[1]+tmp[4590]*kernel[2]+tmp[4688]*kernel[3]+tmp[4689]*kernel[4]+tmp[4690]*kernel[5]+tmp[4788]*kernel[6]+tmp[4789]*kernel[7]+tmp[4790]*kernel[8];
				ans[4690]<=tmp[4589]*kernel[0]+tmp[4590]*kernel[1]+tmp[4591]*kernel[2]+tmp[4689]*kernel[3]+tmp[4690]*kernel[4]+tmp[4691]*kernel[5]+tmp[4789]*kernel[6]+tmp[4790]*kernel[7]+tmp[4791]*kernel[8];
				ans[4691]<=tmp[4590]*kernel[0]+tmp[4591]*kernel[1]+tmp[4592]*kernel[2]+tmp[4690]*kernel[3]+tmp[4691]*kernel[4]+tmp[4692]*kernel[5]+tmp[4790]*kernel[6]+tmp[4791]*kernel[7]+tmp[4792]*kernel[8];
				ans[4692]<=tmp[4591]*kernel[0]+tmp[4592]*kernel[1]+tmp[4593]*kernel[2]+tmp[4691]*kernel[3]+tmp[4692]*kernel[4]+tmp[4693]*kernel[5]+tmp[4791]*kernel[6]+tmp[4792]*kernel[7]+tmp[4793]*kernel[8];
				ans[4693]<=tmp[4592]*kernel[0]+tmp[4593]*kernel[1]+tmp[4594]*kernel[2]+tmp[4692]*kernel[3]+tmp[4693]*kernel[4]+tmp[4694]*kernel[5]+tmp[4792]*kernel[6]+tmp[4793]*kernel[7]+tmp[4794]*kernel[8];
				ans[4694]<=tmp[4593]*kernel[0]+tmp[4594]*kernel[1]+tmp[4595]*kernel[2]+tmp[4693]*kernel[3]+tmp[4694]*kernel[4]+tmp[4695]*kernel[5]+tmp[4793]*kernel[6]+tmp[4794]*kernel[7]+tmp[4795]*kernel[8];
				ans[4695]<=tmp[4594]*kernel[0]+tmp[4595]*kernel[1]+tmp[4596]*kernel[2]+tmp[4694]*kernel[3]+tmp[4695]*kernel[4]+tmp[4696]*kernel[5]+tmp[4794]*kernel[6]+tmp[4795]*kernel[7]+tmp[4796]*kernel[8];
				ans[4696]<=tmp[4595]*kernel[0]+tmp[4596]*kernel[1]+tmp[4597]*kernel[2]+tmp[4695]*kernel[3]+tmp[4696]*kernel[4]+tmp[4697]*kernel[5]+tmp[4795]*kernel[6]+tmp[4796]*kernel[7]+tmp[4797]*kernel[8];
				ans[4697]<=tmp[4596]*kernel[0]+tmp[4597]*kernel[1]+tmp[4598]*kernel[2]+tmp[4696]*kernel[3]+tmp[4697]*kernel[4]+tmp[4698]*kernel[5]+tmp[4796]*kernel[6]+tmp[4797]*kernel[7]+tmp[4798]*kernel[8];
				ans[4698]<=tmp[4597]*kernel[0]+tmp[4598]*kernel[1]+tmp[4599]*kernel[2]+tmp[4697]*kernel[3]+tmp[4698]*kernel[4]+tmp[4699]*kernel[5]+tmp[4797]*kernel[6]+tmp[4798]*kernel[7]+tmp[4799]*kernel[8];
				ans[4699]<=tmp[4598]*kernel[0]+tmp[4599]*kernel[1]+tmp[4698]*kernel[3]+tmp[4699]*kernel[4]+tmp[4798]*kernel[6]+tmp[4799]*kernel[7];
				ans[4700]<=tmp[4600]*kernel[1]+tmp[4601]*kernel[2]+tmp[4700]*kernel[4]+tmp[4701]*kernel[5]+tmp[4800]*kernel[7]+tmp[4801]*kernel[8];
				ans[4701]<=tmp[4600]*kernel[0]+tmp[4601]*kernel[1]+tmp[4602]*kernel[2]+tmp[4700]*kernel[3]+tmp[4701]*kernel[4]+tmp[4702]*kernel[5]+tmp[4800]*kernel[6]+tmp[4801]*kernel[7]+tmp[4802]*kernel[8];
				ans[4702]<=tmp[4601]*kernel[0]+tmp[4602]*kernel[1]+tmp[4603]*kernel[2]+tmp[4701]*kernel[3]+tmp[4702]*kernel[4]+tmp[4703]*kernel[5]+tmp[4801]*kernel[6]+tmp[4802]*kernel[7]+tmp[4803]*kernel[8];
				ans[4703]<=tmp[4602]*kernel[0]+tmp[4603]*kernel[1]+tmp[4604]*kernel[2]+tmp[4702]*kernel[3]+tmp[4703]*kernel[4]+tmp[4704]*kernel[5]+tmp[4802]*kernel[6]+tmp[4803]*kernel[7]+tmp[4804]*kernel[8];
				ans[4704]<=tmp[4603]*kernel[0]+tmp[4604]*kernel[1]+tmp[4605]*kernel[2]+tmp[4703]*kernel[3]+tmp[4704]*kernel[4]+tmp[4705]*kernel[5]+tmp[4803]*kernel[6]+tmp[4804]*kernel[7]+tmp[4805]*kernel[8];
				ans[4705]<=tmp[4604]*kernel[0]+tmp[4605]*kernel[1]+tmp[4606]*kernel[2]+tmp[4704]*kernel[3]+tmp[4705]*kernel[4]+tmp[4706]*kernel[5]+tmp[4804]*kernel[6]+tmp[4805]*kernel[7]+tmp[4806]*kernel[8];
				ans[4706]<=tmp[4605]*kernel[0]+tmp[4606]*kernel[1]+tmp[4607]*kernel[2]+tmp[4705]*kernel[3]+tmp[4706]*kernel[4]+tmp[4707]*kernel[5]+tmp[4805]*kernel[6]+tmp[4806]*kernel[7]+tmp[4807]*kernel[8];
				ans[4707]<=tmp[4606]*kernel[0]+tmp[4607]*kernel[1]+tmp[4608]*kernel[2]+tmp[4706]*kernel[3]+tmp[4707]*kernel[4]+tmp[4708]*kernel[5]+tmp[4806]*kernel[6]+tmp[4807]*kernel[7]+tmp[4808]*kernel[8];
				ans[4708]<=tmp[4607]*kernel[0]+tmp[4608]*kernel[1]+tmp[4609]*kernel[2]+tmp[4707]*kernel[3]+tmp[4708]*kernel[4]+tmp[4709]*kernel[5]+tmp[4807]*kernel[6]+tmp[4808]*kernel[7]+tmp[4809]*kernel[8];
				ans[4709]<=tmp[4608]*kernel[0]+tmp[4609]*kernel[1]+tmp[4610]*kernel[2]+tmp[4708]*kernel[3]+tmp[4709]*kernel[4]+tmp[4710]*kernel[5]+tmp[4808]*kernel[6]+tmp[4809]*kernel[7]+tmp[4810]*kernel[8];
				ans[4710]<=tmp[4609]*kernel[0]+tmp[4610]*kernel[1]+tmp[4611]*kernel[2]+tmp[4709]*kernel[3]+tmp[4710]*kernel[4]+tmp[4711]*kernel[5]+tmp[4809]*kernel[6]+tmp[4810]*kernel[7]+tmp[4811]*kernel[8];
				ans[4711]<=tmp[4610]*kernel[0]+tmp[4611]*kernel[1]+tmp[4612]*kernel[2]+tmp[4710]*kernel[3]+tmp[4711]*kernel[4]+tmp[4712]*kernel[5]+tmp[4810]*kernel[6]+tmp[4811]*kernel[7]+tmp[4812]*kernel[8];
				ans[4712]<=tmp[4611]*kernel[0]+tmp[4612]*kernel[1]+tmp[4613]*kernel[2]+tmp[4711]*kernel[3]+tmp[4712]*kernel[4]+tmp[4713]*kernel[5]+tmp[4811]*kernel[6]+tmp[4812]*kernel[7]+tmp[4813]*kernel[8];
				ans[4713]<=tmp[4612]*kernel[0]+tmp[4613]*kernel[1]+tmp[4614]*kernel[2]+tmp[4712]*kernel[3]+tmp[4713]*kernel[4]+tmp[4714]*kernel[5]+tmp[4812]*kernel[6]+tmp[4813]*kernel[7]+tmp[4814]*kernel[8];
				ans[4714]<=tmp[4613]*kernel[0]+tmp[4614]*kernel[1]+tmp[4615]*kernel[2]+tmp[4713]*kernel[3]+tmp[4714]*kernel[4]+tmp[4715]*kernel[5]+tmp[4813]*kernel[6]+tmp[4814]*kernel[7]+tmp[4815]*kernel[8];
				ans[4715]<=tmp[4614]*kernel[0]+tmp[4615]*kernel[1]+tmp[4616]*kernel[2]+tmp[4714]*kernel[3]+tmp[4715]*kernel[4]+tmp[4716]*kernel[5]+tmp[4814]*kernel[6]+tmp[4815]*kernel[7]+tmp[4816]*kernel[8];
				ans[4716]<=tmp[4615]*kernel[0]+tmp[4616]*kernel[1]+tmp[4617]*kernel[2]+tmp[4715]*kernel[3]+tmp[4716]*kernel[4]+tmp[4717]*kernel[5]+tmp[4815]*kernel[6]+tmp[4816]*kernel[7]+tmp[4817]*kernel[8];
				ans[4717]<=tmp[4616]*kernel[0]+tmp[4617]*kernel[1]+tmp[4618]*kernel[2]+tmp[4716]*kernel[3]+tmp[4717]*kernel[4]+tmp[4718]*kernel[5]+tmp[4816]*kernel[6]+tmp[4817]*kernel[7]+tmp[4818]*kernel[8];
				ans[4718]<=tmp[4617]*kernel[0]+tmp[4618]*kernel[1]+tmp[4619]*kernel[2]+tmp[4717]*kernel[3]+tmp[4718]*kernel[4]+tmp[4719]*kernel[5]+tmp[4817]*kernel[6]+tmp[4818]*kernel[7]+tmp[4819]*kernel[8];
				ans[4719]<=tmp[4618]*kernel[0]+tmp[4619]*kernel[1]+tmp[4620]*kernel[2]+tmp[4718]*kernel[3]+tmp[4719]*kernel[4]+tmp[4720]*kernel[5]+tmp[4818]*kernel[6]+tmp[4819]*kernel[7]+tmp[4820]*kernel[8];
				ans[4720]<=tmp[4619]*kernel[0]+tmp[4620]*kernel[1]+tmp[4621]*kernel[2]+tmp[4719]*kernel[3]+tmp[4720]*kernel[4]+tmp[4721]*kernel[5]+tmp[4819]*kernel[6]+tmp[4820]*kernel[7]+tmp[4821]*kernel[8];
				ans[4721]<=tmp[4620]*kernel[0]+tmp[4621]*kernel[1]+tmp[4622]*kernel[2]+tmp[4720]*kernel[3]+tmp[4721]*kernel[4]+tmp[4722]*kernel[5]+tmp[4820]*kernel[6]+tmp[4821]*kernel[7]+tmp[4822]*kernel[8];
				ans[4722]<=tmp[4621]*kernel[0]+tmp[4622]*kernel[1]+tmp[4623]*kernel[2]+tmp[4721]*kernel[3]+tmp[4722]*kernel[4]+tmp[4723]*kernel[5]+tmp[4821]*kernel[6]+tmp[4822]*kernel[7]+tmp[4823]*kernel[8];
				ans[4723]<=tmp[4622]*kernel[0]+tmp[4623]*kernel[1]+tmp[4624]*kernel[2]+tmp[4722]*kernel[3]+tmp[4723]*kernel[4]+tmp[4724]*kernel[5]+tmp[4822]*kernel[6]+tmp[4823]*kernel[7]+tmp[4824]*kernel[8];
				ans[4724]<=tmp[4623]*kernel[0]+tmp[4624]*kernel[1]+tmp[4625]*kernel[2]+tmp[4723]*kernel[3]+tmp[4724]*kernel[4]+tmp[4725]*kernel[5]+tmp[4823]*kernel[6]+tmp[4824]*kernel[7]+tmp[4825]*kernel[8];
				ans[4725]<=tmp[4624]*kernel[0]+tmp[4625]*kernel[1]+tmp[4626]*kernel[2]+tmp[4724]*kernel[3]+tmp[4725]*kernel[4]+tmp[4726]*kernel[5]+tmp[4824]*kernel[6]+tmp[4825]*kernel[7]+tmp[4826]*kernel[8];
				ans[4726]<=tmp[4625]*kernel[0]+tmp[4626]*kernel[1]+tmp[4627]*kernel[2]+tmp[4725]*kernel[3]+tmp[4726]*kernel[4]+tmp[4727]*kernel[5]+tmp[4825]*kernel[6]+tmp[4826]*kernel[7]+tmp[4827]*kernel[8];
				ans[4727]<=tmp[4626]*kernel[0]+tmp[4627]*kernel[1]+tmp[4628]*kernel[2]+tmp[4726]*kernel[3]+tmp[4727]*kernel[4]+tmp[4728]*kernel[5]+tmp[4826]*kernel[6]+tmp[4827]*kernel[7]+tmp[4828]*kernel[8];
				ans[4728]<=tmp[4627]*kernel[0]+tmp[4628]*kernel[1]+tmp[4629]*kernel[2]+tmp[4727]*kernel[3]+tmp[4728]*kernel[4]+tmp[4729]*kernel[5]+tmp[4827]*kernel[6]+tmp[4828]*kernel[7]+tmp[4829]*kernel[8];
				ans[4729]<=tmp[4628]*kernel[0]+tmp[4629]*kernel[1]+tmp[4630]*kernel[2]+tmp[4728]*kernel[3]+tmp[4729]*kernel[4]+tmp[4730]*kernel[5]+tmp[4828]*kernel[6]+tmp[4829]*kernel[7]+tmp[4830]*kernel[8];
				ans[4730]<=tmp[4629]*kernel[0]+tmp[4630]*kernel[1]+tmp[4631]*kernel[2]+tmp[4729]*kernel[3]+tmp[4730]*kernel[4]+tmp[4731]*kernel[5]+tmp[4829]*kernel[6]+tmp[4830]*kernel[7]+tmp[4831]*kernel[8];
				ans[4731]<=tmp[4630]*kernel[0]+tmp[4631]*kernel[1]+tmp[4632]*kernel[2]+tmp[4730]*kernel[3]+tmp[4731]*kernel[4]+tmp[4732]*kernel[5]+tmp[4830]*kernel[6]+tmp[4831]*kernel[7]+tmp[4832]*kernel[8];
				ans[4732]<=tmp[4631]*kernel[0]+tmp[4632]*kernel[1]+tmp[4633]*kernel[2]+tmp[4731]*kernel[3]+tmp[4732]*kernel[4]+tmp[4733]*kernel[5]+tmp[4831]*kernel[6]+tmp[4832]*kernel[7]+tmp[4833]*kernel[8];
				ans[4733]<=tmp[4632]*kernel[0]+tmp[4633]*kernel[1]+tmp[4634]*kernel[2]+tmp[4732]*kernel[3]+tmp[4733]*kernel[4]+tmp[4734]*kernel[5]+tmp[4832]*kernel[6]+tmp[4833]*kernel[7]+tmp[4834]*kernel[8];
				ans[4734]<=tmp[4633]*kernel[0]+tmp[4634]*kernel[1]+tmp[4635]*kernel[2]+tmp[4733]*kernel[3]+tmp[4734]*kernel[4]+tmp[4735]*kernel[5]+tmp[4833]*kernel[6]+tmp[4834]*kernel[7]+tmp[4835]*kernel[8];
				ans[4735]<=tmp[4634]*kernel[0]+tmp[4635]*kernel[1]+tmp[4636]*kernel[2]+tmp[4734]*kernel[3]+tmp[4735]*kernel[4]+tmp[4736]*kernel[5]+tmp[4834]*kernel[6]+tmp[4835]*kernel[7]+tmp[4836]*kernel[8];
				ans[4736]<=tmp[4635]*kernel[0]+tmp[4636]*kernel[1]+tmp[4637]*kernel[2]+tmp[4735]*kernel[3]+tmp[4736]*kernel[4]+tmp[4737]*kernel[5]+tmp[4835]*kernel[6]+tmp[4836]*kernel[7]+tmp[4837]*kernel[8];
				ans[4737]<=tmp[4636]*kernel[0]+tmp[4637]*kernel[1]+tmp[4638]*kernel[2]+tmp[4736]*kernel[3]+tmp[4737]*kernel[4]+tmp[4738]*kernel[5]+tmp[4836]*kernel[6]+tmp[4837]*kernel[7]+tmp[4838]*kernel[8];
				ans[4738]<=tmp[4637]*kernel[0]+tmp[4638]*kernel[1]+tmp[4639]*kernel[2]+tmp[4737]*kernel[3]+tmp[4738]*kernel[4]+tmp[4739]*kernel[5]+tmp[4837]*kernel[6]+tmp[4838]*kernel[7]+tmp[4839]*kernel[8];
				ans[4739]<=tmp[4638]*kernel[0]+tmp[4639]*kernel[1]+tmp[4640]*kernel[2]+tmp[4738]*kernel[3]+tmp[4739]*kernel[4]+tmp[4740]*kernel[5]+tmp[4838]*kernel[6]+tmp[4839]*kernel[7]+tmp[4840]*kernel[8];
				ans[4740]<=tmp[4639]*kernel[0]+tmp[4640]*kernel[1]+tmp[4641]*kernel[2]+tmp[4739]*kernel[3]+tmp[4740]*kernel[4]+tmp[4741]*kernel[5]+tmp[4839]*kernel[6]+tmp[4840]*kernel[7]+tmp[4841]*kernel[8];
				ans[4741]<=tmp[4640]*kernel[0]+tmp[4641]*kernel[1]+tmp[4642]*kernel[2]+tmp[4740]*kernel[3]+tmp[4741]*kernel[4]+tmp[4742]*kernel[5]+tmp[4840]*kernel[6]+tmp[4841]*kernel[7]+tmp[4842]*kernel[8];
				ans[4742]<=tmp[4641]*kernel[0]+tmp[4642]*kernel[1]+tmp[4643]*kernel[2]+tmp[4741]*kernel[3]+tmp[4742]*kernel[4]+tmp[4743]*kernel[5]+tmp[4841]*kernel[6]+tmp[4842]*kernel[7]+tmp[4843]*kernel[8];
				ans[4743]<=tmp[4642]*kernel[0]+tmp[4643]*kernel[1]+tmp[4644]*kernel[2]+tmp[4742]*kernel[3]+tmp[4743]*kernel[4]+tmp[4744]*kernel[5]+tmp[4842]*kernel[6]+tmp[4843]*kernel[7]+tmp[4844]*kernel[8];
				ans[4744]<=tmp[4643]*kernel[0]+tmp[4644]*kernel[1]+tmp[4645]*kernel[2]+tmp[4743]*kernel[3]+tmp[4744]*kernel[4]+tmp[4745]*kernel[5]+tmp[4843]*kernel[6]+tmp[4844]*kernel[7]+tmp[4845]*kernel[8];
				ans[4745]<=tmp[4644]*kernel[0]+tmp[4645]*kernel[1]+tmp[4646]*kernel[2]+tmp[4744]*kernel[3]+tmp[4745]*kernel[4]+tmp[4746]*kernel[5]+tmp[4844]*kernel[6]+tmp[4845]*kernel[7]+tmp[4846]*kernel[8];
				ans[4746]<=tmp[4645]*kernel[0]+tmp[4646]*kernel[1]+tmp[4647]*kernel[2]+tmp[4745]*kernel[3]+tmp[4746]*kernel[4]+tmp[4747]*kernel[5]+tmp[4845]*kernel[6]+tmp[4846]*kernel[7]+tmp[4847]*kernel[8];
				ans[4747]<=tmp[4646]*kernel[0]+tmp[4647]*kernel[1]+tmp[4648]*kernel[2]+tmp[4746]*kernel[3]+tmp[4747]*kernel[4]+tmp[4748]*kernel[5]+tmp[4846]*kernel[6]+tmp[4847]*kernel[7]+tmp[4848]*kernel[8];
				ans[4748]<=tmp[4647]*kernel[0]+tmp[4648]*kernel[1]+tmp[4649]*kernel[2]+tmp[4747]*kernel[3]+tmp[4748]*kernel[4]+tmp[4749]*kernel[5]+tmp[4847]*kernel[6]+tmp[4848]*kernel[7]+tmp[4849]*kernel[8];
				ans[4749]<=tmp[4648]*kernel[0]+tmp[4649]*kernel[1]+tmp[4650]*kernel[2]+tmp[4748]*kernel[3]+tmp[4749]*kernel[4]+tmp[4750]*kernel[5]+tmp[4848]*kernel[6]+tmp[4849]*kernel[7]+tmp[4850]*kernel[8];
				ans[4750]<=tmp[4649]*kernel[0]+tmp[4650]*kernel[1]+tmp[4651]*kernel[2]+tmp[4749]*kernel[3]+tmp[4750]*kernel[4]+tmp[4751]*kernel[5]+tmp[4849]*kernel[6]+tmp[4850]*kernel[7]+tmp[4851]*kernel[8];
				ans[4751]<=tmp[4650]*kernel[0]+tmp[4651]*kernel[1]+tmp[4652]*kernel[2]+tmp[4750]*kernel[3]+tmp[4751]*kernel[4]+tmp[4752]*kernel[5]+tmp[4850]*kernel[6]+tmp[4851]*kernel[7]+tmp[4852]*kernel[8];
				ans[4752]<=tmp[4651]*kernel[0]+tmp[4652]*kernel[1]+tmp[4653]*kernel[2]+tmp[4751]*kernel[3]+tmp[4752]*kernel[4]+tmp[4753]*kernel[5]+tmp[4851]*kernel[6]+tmp[4852]*kernel[7]+tmp[4853]*kernel[8];
				ans[4753]<=tmp[4652]*kernel[0]+tmp[4653]*kernel[1]+tmp[4654]*kernel[2]+tmp[4752]*kernel[3]+tmp[4753]*kernel[4]+tmp[4754]*kernel[5]+tmp[4852]*kernel[6]+tmp[4853]*kernel[7]+tmp[4854]*kernel[8];
				ans[4754]<=tmp[4653]*kernel[0]+tmp[4654]*kernel[1]+tmp[4655]*kernel[2]+tmp[4753]*kernel[3]+tmp[4754]*kernel[4]+tmp[4755]*kernel[5]+tmp[4853]*kernel[6]+tmp[4854]*kernel[7]+tmp[4855]*kernel[8];
				ans[4755]<=tmp[4654]*kernel[0]+tmp[4655]*kernel[1]+tmp[4656]*kernel[2]+tmp[4754]*kernel[3]+tmp[4755]*kernel[4]+tmp[4756]*kernel[5]+tmp[4854]*kernel[6]+tmp[4855]*kernel[7]+tmp[4856]*kernel[8];
				ans[4756]<=tmp[4655]*kernel[0]+tmp[4656]*kernel[1]+tmp[4657]*kernel[2]+tmp[4755]*kernel[3]+tmp[4756]*kernel[4]+tmp[4757]*kernel[5]+tmp[4855]*kernel[6]+tmp[4856]*kernel[7]+tmp[4857]*kernel[8];
				ans[4757]<=tmp[4656]*kernel[0]+tmp[4657]*kernel[1]+tmp[4658]*kernel[2]+tmp[4756]*kernel[3]+tmp[4757]*kernel[4]+tmp[4758]*kernel[5]+tmp[4856]*kernel[6]+tmp[4857]*kernel[7]+tmp[4858]*kernel[8];
				ans[4758]<=tmp[4657]*kernel[0]+tmp[4658]*kernel[1]+tmp[4659]*kernel[2]+tmp[4757]*kernel[3]+tmp[4758]*kernel[4]+tmp[4759]*kernel[5]+tmp[4857]*kernel[6]+tmp[4858]*kernel[7]+tmp[4859]*kernel[8];
				ans[4759]<=tmp[4658]*kernel[0]+tmp[4659]*kernel[1]+tmp[4660]*kernel[2]+tmp[4758]*kernel[3]+tmp[4759]*kernel[4]+tmp[4760]*kernel[5]+tmp[4858]*kernel[6]+tmp[4859]*kernel[7]+tmp[4860]*kernel[8];
				ans[4760]<=tmp[4659]*kernel[0]+tmp[4660]*kernel[1]+tmp[4661]*kernel[2]+tmp[4759]*kernel[3]+tmp[4760]*kernel[4]+tmp[4761]*kernel[5]+tmp[4859]*kernel[6]+tmp[4860]*kernel[7]+tmp[4861]*kernel[8];
				ans[4761]<=tmp[4660]*kernel[0]+tmp[4661]*kernel[1]+tmp[4662]*kernel[2]+tmp[4760]*kernel[3]+tmp[4761]*kernel[4]+tmp[4762]*kernel[5]+tmp[4860]*kernel[6]+tmp[4861]*kernel[7]+tmp[4862]*kernel[8];
				ans[4762]<=tmp[4661]*kernel[0]+tmp[4662]*kernel[1]+tmp[4663]*kernel[2]+tmp[4761]*kernel[3]+tmp[4762]*kernel[4]+tmp[4763]*kernel[5]+tmp[4861]*kernel[6]+tmp[4862]*kernel[7]+tmp[4863]*kernel[8];
				ans[4763]<=tmp[4662]*kernel[0]+tmp[4663]*kernel[1]+tmp[4664]*kernel[2]+tmp[4762]*kernel[3]+tmp[4763]*kernel[4]+tmp[4764]*kernel[5]+tmp[4862]*kernel[6]+tmp[4863]*kernel[7]+tmp[4864]*kernel[8];
				ans[4764]<=tmp[4663]*kernel[0]+tmp[4664]*kernel[1]+tmp[4665]*kernel[2]+tmp[4763]*kernel[3]+tmp[4764]*kernel[4]+tmp[4765]*kernel[5]+tmp[4863]*kernel[6]+tmp[4864]*kernel[7]+tmp[4865]*kernel[8];
				ans[4765]<=tmp[4664]*kernel[0]+tmp[4665]*kernel[1]+tmp[4666]*kernel[2]+tmp[4764]*kernel[3]+tmp[4765]*kernel[4]+tmp[4766]*kernel[5]+tmp[4864]*kernel[6]+tmp[4865]*kernel[7]+tmp[4866]*kernel[8];
				ans[4766]<=tmp[4665]*kernel[0]+tmp[4666]*kernel[1]+tmp[4667]*kernel[2]+tmp[4765]*kernel[3]+tmp[4766]*kernel[4]+tmp[4767]*kernel[5]+tmp[4865]*kernel[6]+tmp[4866]*kernel[7]+tmp[4867]*kernel[8];
				ans[4767]<=tmp[4666]*kernel[0]+tmp[4667]*kernel[1]+tmp[4668]*kernel[2]+tmp[4766]*kernel[3]+tmp[4767]*kernel[4]+tmp[4768]*kernel[5]+tmp[4866]*kernel[6]+tmp[4867]*kernel[7]+tmp[4868]*kernel[8];
				ans[4768]<=tmp[4667]*kernel[0]+tmp[4668]*kernel[1]+tmp[4669]*kernel[2]+tmp[4767]*kernel[3]+tmp[4768]*kernel[4]+tmp[4769]*kernel[5]+tmp[4867]*kernel[6]+tmp[4868]*kernel[7]+tmp[4869]*kernel[8];
				ans[4769]<=tmp[4668]*kernel[0]+tmp[4669]*kernel[1]+tmp[4670]*kernel[2]+tmp[4768]*kernel[3]+tmp[4769]*kernel[4]+tmp[4770]*kernel[5]+tmp[4868]*kernel[6]+tmp[4869]*kernel[7]+tmp[4870]*kernel[8];
				ans[4770]<=tmp[4669]*kernel[0]+tmp[4670]*kernel[1]+tmp[4671]*kernel[2]+tmp[4769]*kernel[3]+tmp[4770]*kernel[4]+tmp[4771]*kernel[5]+tmp[4869]*kernel[6]+tmp[4870]*kernel[7]+tmp[4871]*kernel[8];
				ans[4771]<=tmp[4670]*kernel[0]+tmp[4671]*kernel[1]+tmp[4672]*kernel[2]+tmp[4770]*kernel[3]+tmp[4771]*kernel[4]+tmp[4772]*kernel[5]+tmp[4870]*kernel[6]+tmp[4871]*kernel[7]+tmp[4872]*kernel[8];
				ans[4772]<=tmp[4671]*kernel[0]+tmp[4672]*kernel[1]+tmp[4673]*kernel[2]+tmp[4771]*kernel[3]+tmp[4772]*kernel[4]+tmp[4773]*kernel[5]+tmp[4871]*kernel[6]+tmp[4872]*kernel[7]+tmp[4873]*kernel[8];
				ans[4773]<=tmp[4672]*kernel[0]+tmp[4673]*kernel[1]+tmp[4674]*kernel[2]+tmp[4772]*kernel[3]+tmp[4773]*kernel[4]+tmp[4774]*kernel[5]+tmp[4872]*kernel[6]+tmp[4873]*kernel[7]+tmp[4874]*kernel[8];
				ans[4774]<=tmp[4673]*kernel[0]+tmp[4674]*kernel[1]+tmp[4675]*kernel[2]+tmp[4773]*kernel[3]+tmp[4774]*kernel[4]+tmp[4775]*kernel[5]+tmp[4873]*kernel[6]+tmp[4874]*kernel[7]+tmp[4875]*kernel[8];
				ans[4775]<=tmp[4674]*kernel[0]+tmp[4675]*kernel[1]+tmp[4676]*kernel[2]+tmp[4774]*kernel[3]+tmp[4775]*kernel[4]+tmp[4776]*kernel[5]+tmp[4874]*kernel[6]+tmp[4875]*kernel[7]+tmp[4876]*kernel[8];
				ans[4776]<=tmp[4675]*kernel[0]+tmp[4676]*kernel[1]+tmp[4677]*kernel[2]+tmp[4775]*kernel[3]+tmp[4776]*kernel[4]+tmp[4777]*kernel[5]+tmp[4875]*kernel[6]+tmp[4876]*kernel[7]+tmp[4877]*kernel[8];
				ans[4777]<=tmp[4676]*kernel[0]+tmp[4677]*kernel[1]+tmp[4678]*kernel[2]+tmp[4776]*kernel[3]+tmp[4777]*kernel[4]+tmp[4778]*kernel[5]+tmp[4876]*kernel[6]+tmp[4877]*kernel[7]+tmp[4878]*kernel[8];
				ans[4778]<=tmp[4677]*kernel[0]+tmp[4678]*kernel[1]+tmp[4679]*kernel[2]+tmp[4777]*kernel[3]+tmp[4778]*kernel[4]+tmp[4779]*kernel[5]+tmp[4877]*kernel[6]+tmp[4878]*kernel[7]+tmp[4879]*kernel[8];
				ans[4779]<=tmp[4678]*kernel[0]+tmp[4679]*kernel[1]+tmp[4680]*kernel[2]+tmp[4778]*kernel[3]+tmp[4779]*kernel[4]+tmp[4780]*kernel[5]+tmp[4878]*kernel[6]+tmp[4879]*kernel[7]+tmp[4880]*kernel[8];
				ans[4780]<=tmp[4679]*kernel[0]+tmp[4680]*kernel[1]+tmp[4681]*kernel[2]+tmp[4779]*kernel[3]+tmp[4780]*kernel[4]+tmp[4781]*kernel[5]+tmp[4879]*kernel[6]+tmp[4880]*kernel[7]+tmp[4881]*kernel[8];
				ans[4781]<=tmp[4680]*kernel[0]+tmp[4681]*kernel[1]+tmp[4682]*kernel[2]+tmp[4780]*kernel[3]+tmp[4781]*kernel[4]+tmp[4782]*kernel[5]+tmp[4880]*kernel[6]+tmp[4881]*kernel[7]+tmp[4882]*kernel[8];
				ans[4782]<=tmp[4681]*kernel[0]+tmp[4682]*kernel[1]+tmp[4683]*kernel[2]+tmp[4781]*kernel[3]+tmp[4782]*kernel[4]+tmp[4783]*kernel[5]+tmp[4881]*kernel[6]+tmp[4882]*kernel[7]+tmp[4883]*kernel[8];
				ans[4783]<=tmp[4682]*kernel[0]+tmp[4683]*kernel[1]+tmp[4684]*kernel[2]+tmp[4782]*kernel[3]+tmp[4783]*kernel[4]+tmp[4784]*kernel[5]+tmp[4882]*kernel[6]+tmp[4883]*kernel[7]+tmp[4884]*kernel[8];
				ans[4784]<=tmp[4683]*kernel[0]+tmp[4684]*kernel[1]+tmp[4685]*kernel[2]+tmp[4783]*kernel[3]+tmp[4784]*kernel[4]+tmp[4785]*kernel[5]+tmp[4883]*kernel[6]+tmp[4884]*kernel[7]+tmp[4885]*kernel[8];
				ans[4785]<=tmp[4684]*kernel[0]+tmp[4685]*kernel[1]+tmp[4686]*kernel[2]+tmp[4784]*kernel[3]+tmp[4785]*kernel[4]+tmp[4786]*kernel[5]+tmp[4884]*kernel[6]+tmp[4885]*kernel[7]+tmp[4886]*kernel[8];
				ans[4786]<=tmp[4685]*kernel[0]+tmp[4686]*kernel[1]+tmp[4687]*kernel[2]+tmp[4785]*kernel[3]+tmp[4786]*kernel[4]+tmp[4787]*kernel[5]+tmp[4885]*kernel[6]+tmp[4886]*kernel[7]+tmp[4887]*kernel[8];
				ans[4787]<=tmp[4686]*kernel[0]+tmp[4687]*kernel[1]+tmp[4688]*kernel[2]+tmp[4786]*kernel[3]+tmp[4787]*kernel[4]+tmp[4788]*kernel[5]+tmp[4886]*kernel[6]+tmp[4887]*kernel[7]+tmp[4888]*kernel[8];
				ans[4788]<=tmp[4687]*kernel[0]+tmp[4688]*kernel[1]+tmp[4689]*kernel[2]+tmp[4787]*kernel[3]+tmp[4788]*kernel[4]+tmp[4789]*kernel[5]+tmp[4887]*kernel[6]+tmp[4888]*kernel[7]+tmp[4889]*kernel[8];
				ans[4789]<=tmp[4688]*kernel[0]+tmp[4689]*kernel[1]+tmp[4690]*kernel[2]+tmp[4788]*kernel[3]+tmp[4789]*kernel[4]+tmp[4790]*kernel[5]+tmp[4888]*kernel[6]+tmp[4889]*kernel[7]+tmp[4890]*kernel[8];
				ans[4790]<=tmp[4689]*kernel[0]+tmp[4690]*kernel[1]+tmp[4691]*kernel[2]+tmp[4789]*kernel[3]+tmp[4790]*kernel[4]+tmp[4791]*kernel[5]+tmp[4889]*kernel[6]+tmp[4890]*kernel[7]+tmp[4891]*kernel[8];
				ans[4791]<=tmp[4690]*kernel[0]+tmp[4691]*kernel[1]+tmp[4692]*kernel[2]+tmp[4790]*kernel[3]+tmp[4791]*kernel[4]+tmp[4792]*kernel[5]+tmp[4890]*kernel[6]+tmp[4891]*kernel[7]+tmp[4892]*kernel[8];
				ans[4792]<=tmp[4691]*kernel[0]+tmp[4692]*kernel[1]+tmp[4693]*kernel[2]+tmp[4791]*kernel[3]+tmp[4792]*kernel[4]+tmp[4793]*kernel[5]+tmp[4891]*kernel[6]+tmp[4892]*kernel[7]+tmp[4893]*kernel[8];
				ans[4793]<=tmp[4692]*kernel[0]+tmp[4693]*kernel[1]+tmp[4694]*kernel[2]+tmp[4792]*kernel[3]+tmp[4793]*kernel[4]+tmp[4794]*kernel[5]+tmp[4892]*kernel[6]+tmp[4893]*kernel[7]+tmp[4894]*kernel[8];
				ans[4794]<=tmp[4693]*kernel[0]+tmp[4694]*kernel[1]+tmp[4695]*kernel[2]+tmp[4793]*kernel[3]+tmp[4794]*kernel[4]+tmp[4795]*kernel[5]+tmp[4893]*kernel[6]+tmp[4894]*kernel[7]+tmp[4895]*kernel[8];
				ans[4795]<=tmp[4694]*kernel[0]+tmp[4695]*kernel[1]+tmp[4696]*kernel[2]+tmp[4794]*kernel[3]+tmp[4795]*kernel[4]+tmp[4796]*kernel[5]+tmp[4894]*kernel[6]+tmp[4895]*kernel[7]+tmp[4896]*kernel[8];
				ans[4796]<=tmp[4695]*kernel[0]+tmp[4696]*kernel[1]+tmp[4697]*kernel[2]+tmp[4795]*kernel[3]+tmp[4796]*kernel[4]+tmp[4797]*kernel[5]+tmp[4895]*kernel[6]+tmp[4896]*kernel[7]+tmp[4897]*kernel[8];
				ans[4797]<=tmp[4696]*kernel[0]+tmp[4697]*kernel[1]+tmp[4698]*kernel[2]+tmp[4796]*kernel[3]+tmp[4797]*kernel[4]+tmp[4798]*kernel[5]+tmp[4896]*kernel[6]+tmp[4897]*kernel[7]+tmp[4898]*kernel[8];
				ans[4798]<=tmp[4697]*kernel[0]+tmp[4698]*kernel[1]+tmp[4699]*kernel[2]+tmp[4797]*kernel[3]+tmp[4798]*kernel[4]+tmp[4799]*kernel[5]+tmp[4897]*kernel[6]+tmp[4898]*kernel[7]+tmp[4899]*kernel[8];
				ans[4799]<=tmp[4698]*kernel[0]+tmp[4699]*kernel[1]+tmp[4798]*kernel[3]+tmp[4799]*kernel[4]+tmp[4898]*kernel[6]+tmp[4899]*kernel[7];
				ans[4800]<=tmp[4700]*kernel[1]+tmp[4701]*kernel[2]+tmp[4800]*kernel[4]+tmp[4801]*kernel[5]+tmp[4900]*kernel[7]+tmp[4901]*kernel[8];
				ans[4801]<=tmp[4700]*kernel[0]+tmp[4701]*kernel[1]+tmp[4702]*kernel[2]+tmp[4800]*kernel[3]+tmp[4801]*kernel[4]+tmp[4802]*kernel[5]+tmp[4900]*kernel[6]+tmp[4901]*kernel[7]+tmp[4902]*kernel[8];
				ans[4802]<=tmp[4701]*kernel[0]+tmp[4702]*kernel[1]+tmp[4703]*kernel[2]+tmp[4801]*kernel[3]+tmp[4802]*kernel[4]+tmp[4803]*kernel[5]+tmp[4901]*kernel[6]+tmp[4902]*kernel[7]+tmp[4903]*kernel[8];
				ans[4803]<=tmp[4702]*kernel[0]+tmp[4703]*kernel[1]+tmp[4704]*kernel[2]+tmp[4802]*kernel[3]+tmp[4803]*kernel[4]+tmp[4804]*kernel[5]+tmp[4902]*kernel[6]+tmp[4903]*kernel[7]+tmp[4904]*kernel[8];
				ans[4804]<=tmp[4703]*kernel[0]+tmp[4704]*kernel[1]+tmp[4705]*kernel[2]+tmp[4803]*kernel[3]+tmp[4804]*kernel[4]+tmp[4805]*kernel[5]+tmp[4903]*kernel[6]+tmp[4904]*kernel[7]+tmp[4905]*kernel[8];
				ans[4805]<=tmp[4704]*kernel[0]+tmp[4705]*kernel[1]+tmp[4706]*kernel[2]+tmp[4804]*kernel[3]+tmp[4805]*kernel[4]+tmp[4806]*kernel[5]+tmp[4904]*kernel[6]+tmp[4905]*kernel[7]+tmp[4906]*kernel[8];
				ans[4806]<=tmp[4705]*kernel[0]+tmp[4706]*kernel[1]+tmp[4707]*kernel[2]+tmp[4805]*kernel[3]+tmp[4806]*kernel[4]+tmp[4807]*kernel[5]+tmp[4905]*kernel[6]+tmp[4906]*kernel[7]+tmp[4907]*kernel[8];
				ans[4807]<=tmp[4706]*kernel[0]+tmp[4707]*kernel[1]+tmp[4708]*kernel[2]+tmp[4806]*kernel[3]+tmp[4807]*kernel[4]+tmp[4808]*kernel[5]+tmp[4906]*kernel[6]+tmp[4907]*kernel[7]+tmp[4908]*kernel[8];
				ans[4808]<=tmp[4707]*kernel[0]+tmp[4708]*kernel[1]+tmp[4709]*kernel[2]+tmp[4807]*kernel[3]+tmp[4808]*kernel[4]+tmp[4809]*kernel[5]+tmp[4907]*kernel[6]+tmp[4908]*kernel[7]+tmp[4909]*kernel[8];
				ans[4809]<=tmp[4708]*kernel[0]+tmp[4709]*kernel[1]+tmp[4710]*kernel[2]+tmp[4808]*kernel[3]+tmp[4809]*kernel[4]+tmp[4810]*kernel[5]+tmp[4908]*kernel[6]+tmp[4909]*kernel[7]+tmp[4910]*kernel[8];
				ans[4810]<=tmp[4709]*kernel[0]+tmp[4710]*kernel[1]+tmp[4711]*kernel[2]+tmp[4809]*kernel[3]+tmp[4810]*kernel[4]+tmp[4811]*kernel[5]+tmp[4909]*kernel[6]+tmp[4910]*kernel[7]+tmp[4911]*kernel[8];
				ans[4811]<=tmp[4710]*kernel[0]+tmp[4711]*kernel[1]+tmp[4712]*kernel[2]+tmp[4810]*kernel[3]+tmp[4811]*kernel[4]+tmp[4812]*kernel[5]+tmp[4910]*kernel[6]+tmp[4911]*kernel[7]+tmp[4912]*kernel[8];
				ans[4812]<=tmp[4711]*kernel[0]+tmp[4712]*kernel[1]+tmp[4713]*kernel[2]+tmp[4811]*kernel[3]+tmp[4812]*kernel[4]+tmp[4813]*kernel[5]+tmp[4911]*kernel[6]+tmp[4912]*kernel[7]+tmp[4913]*kernel[8];
				ans[4813]<=tmp[4712]*kernel[0]+tmp[4713]*kernel[1]+tmp[4714]*kernel[2]+tmp[4812]*kernel[3]+tmp[4813]*kernel[4]+tmp[4814]*kernel[5]+tmp[4912]*kernel[6]+tmp[4913]*kernel[7]+tmp[4914]*kernel[8];
				ans[4814]<=tmp[4713]*kernel[0]+tmp[4714]*kernel[1]+tmp[4715]*kernel[2]+tmp[4813]*kernel[3]+tmp[4814]*kernel[4]+tmp[4815]*kernel[5]+tmp[4913]*kernel[6]+tmp[4914]*kernel[7]+tmp[4915]*kernel[8];
				ans[4815]<=tmp[4714]*kernel[0]+tmp[4715]*kernel[1]+tmp[4716]*kernel[2]+tmp[4814]*kernel[3]+tmp[4815]*kernel[4]+tmp[4816]*kernel[5]+tmp[4914]*kernel[6]+tmp[4915]*kernel[7]+tmp[4916]*kernel[8];
				ans[4816]<=tmp[4715]*kernel[0]+tmp[4716]*kernel[1]+tmp[4717]*kernel[2]+tmp[4815]*kernel[3]+tmp[4816]*kernel[4]+tmp[4817]*kernel[5]+tmp[4915]*kernel[6]+tmp[4916]*kernel[7]+tmp[4917]*kernel[8];
				ans[4817]<=tmp[4716]*kernel[0]+tmp[4717]*kernel[1]+tmp[4718]*kernel[2]+tmp[4816]*kernel[3]+tmp[4817]*kernel[4]+tmp[4818]*kernel[5]+tmp[4916]*kernel[6]+tmp[4917]*kernel[7]+tmp[4918]*kernel[8];
				ans[4818]<=tmp[4717]*kernel[0]+tmp[4718]*kernel[1]+tmp[4719]*kernel[2]+tmp[4817]*kernel[3]+tmp[4818]*kernel[4]+tmp[4819]*kernel[5]+tmp[4917]*kernel[6]+tmp[4918]*kernel[7]+tmp[4919]*kernel[8];
				ans[4819]<=tmp[4718]*kernel[0]+tmp[4719]*kernel[1]+tmp[4720]*kernel[2]+tmp[4818]*kernel[3]+tmp[4819]*kernel[4]+tmp[4820]*kernel[5]+tmp[4918]*kernel[6]+tmp[4919]*kernel[7]+tmp[4920]*kernel[8];
				ans[4820]<=tmp[4719]*kernel[0]+tmp[4720]*kernel[1]+tmp[4721]*kernel[2]+tmp[4819]*kernel[3]+tmp[4820]*kernel[4]+tmp[4821]*kernel[5]+tmp[4919]*kernel[6]+tmp[4920]*kernel[7]+tmp[4921]*kernel[8];
				ans[4821]<=tmp[4720]*kernel[0]+tmp[4721]*kernel[1]+tmp[4722]*kernel[2]+tmp[4820]*kernel[3]+tmp[4821]*kernel[4]+tmp[4822]*kernel[5]+tmp[4920]*kernel[6]+tmp[4921]*kernel[7]+tmp[4922]*kernel[8];
				ans[4822]<=tmp[4721]*kernel[0]+tmp[4722]*kernel[1]+tmp[4723]*kernel[2]+tmp[4821]*kernel[3]+tmp[4822]*kernel[4]+tmp[4823]*kernel[5]+tmp[4921]*kernel[6]+tmp[4922]*kernel[7]+tmp[4923]*kernel[8];
				ans[4823]<=tmp[4722]*kernel[0]+tmp[4723]*kernel[1]+tmp[4724]*kernel[2]+tmp[4822]*kernel[3]+tmp[4823]*kernel[4]+tmp[4824]*kernel[5]+tmp[4922]*kernel[6]+tmp[4923]*kernel[7]+tmp[4924]*kernel[8];
				ans[4824]<=tmp[4723]*kernel[0]+tmp[4724]*kernel[1]+tmp[4725]*kernel[2]+tmp[4823]*kernel[3]+tmp[4824]*kernel[4]+tmp[4825]*kernel[5]+tmp[4923]*kernel[6]+tmp[4924]*kernel[7]+tmp[4925]*kernel[8];
				ans[4825]<=tmp[4724]*kernel[0]+tmp[4725]*kernel[1]+tmp[4726]*kernel[2]+tmp[4824]*kernel[3]+tmp[4825]*kernel[4]+tmp[4826]*kernel[5]+tmp[4924]*kernel[6]+tmp[4925]*kernel[7]+tmp[4926]*kernel[8];
				ans[4826]<=tmp[4725]*kernel[0]+tmp[4726]*kernel[1]+tmp[4727]*kernel[2]+tmp[4825]*kernel[3]+tmp[4826]*kernel[4]+tmp[4827]*kernel[5]+tmp[4925]*kernel[6]+tmp[4926]*kernel[7]+tmp[4927]*kernel[8];
				ans[4827]<=tmp[4726]*kernel[0]+tmp[4727]*kernel[1]+tmp[4728]*kernel[2]+tmp[4826]*kernel[3]+tmp[4827]*kernel[4]+tmp[4828]*kernel[5]+tmp[4926]*kernel[6]+tmp[4927]*kernel[7]+tmp[4928]*kernel[8];
				ans[4828]<=tmp[4727]*kernel[0]+tmp[4728]*kernel[1]+tmp[4729]*kernel[2]+tmp[4827]*kernel[3]+tmp[4828]*kernel[4]+tmp[4829]*kernel[5]+tmp[4927]*kernel[6]+tmp[4928]*kernel[7]+tmp[4929]*kernel[8];
				ans[4829]<=tmp[4728]*kernel[0]+tmp[4729]*kernel[1]+tmp[4730]*kernel[2]+tmp[4828]*kernel[3]+tmp[4829]*kernel[4]+tmp[4830]*kernel[5]+tmp[4928]*kernel[6]+tmp[4929]*kernel[7]+tmp[4930]*kernel[8];
				ans[4830]<=tmp[4729]*kernel[0]+tmp[4730]*kernel[1]+tmp[4731]*kernel[2]+tmp[4829]*kernel[3]+tmp[4830]*kernel[4]+tmp[4831]*kernel[5]+tmp[4929]*kernel[6]+tmp[4930]*kernel[7]+tmp[4931]*kernel[8];
				ans[4831]<=tmp[4730]*kernel[0]+tmp[4731]*kernel[1]+tmp[4732]*kernel[2]+tmp[4830]*kernel[3]+tmp[4831]*kernel[4]+tmp[4832]*kernel[5]+tmp[4930]*kernel[6]+tmp[4931]*kernel[7]+tmp[4932]*kernel[8];
				ans[4832]<=tmp[4731]*kernel[0]+tmp[4732]*kernel[1]+tmp[4733]*kernel[2]+tmp[4831]*kernel[3]+tmp[4832]*kernel[4]+tmp[4833]*kernel[5]+tmp[4931]*kernel[6]+tmp[4932]*kernel[7]+tmp[4933]*kernel[8];
				ans[4833]<=tmp[4732]*kernel[0]+tmp[4733]*kernel[1]+tmp[4734]*kernel[2]+tmp[4832]*kernel[3]+tmp[4833]*kernel[4]+tmp[4834]*kernel[5]+tmp[4932]*kernel[6]+tmp[4933]*kernel[7]+tmp[4934]*kernel[8];
				ans[4834]<=tmp[4733]*kernel[0]+tmp[4734]*kernel[1]+tmp[4735]*kernel[2]+tmp[4833]*kernel[3]+tmp[4834]*kernel[4]+tmp[4835]*kernel[5]+tmp[4933]*kernel[6]+tmp[4934]*kernel[7]+tmp[4935]*kernel[8];
				ans[4835]<=tmp[4734]*kernel[0]+tmp[4735]*kernel[1]+tmp[4736]*kernel[2]+tmp[4834]*kernel[3]+tmp[4835]*kernel[4]+tmp[4836]*kernel[5]+tmp[4934]*kernel[6]+tmp[4935]*kernel[7]+tmp[4936]*kernel[8];
				ans[4836]<=tmp[4735]*kernel[0]+tmp[4736]*kernel[1]+tmp[4737]*kernel[2]+tmp[4835]*kernel[3]+tmp[4836]*kernel[4]+tmp[4837]*kernel[5]+tmp[4935]*kernel[6]+tmp[4936]*kernel[7]+tmp[4937]*kernel[8];
				ans[4837]<=tmp[4736]*kernel[0]+tmp[4737]*kernel[1]+tmp[4738]*kernel[2]+tmp[4836]*kernel[3]+tmp[4837]*kernel[4]+tmp[4838]*kernel[5]+tmp[4936]*kernel[6]+tmp[4937]*kernel[7]+tmp[4938]*kernel[8];
				ans[4838]<=tmp[4737]*kernel[0]+tmp[4738]*kernel[1]+tmp[4739]*kernel[2]+tmp[4837]*kernel[3]+tmp[4838]*kernel[4]+tmp[4839]*kernel[5]+tmp[4937]*kernel[6]+tmp[4938]*kernel[7]+tmp[4939]*kernel[8];
				ans[4839]<=tmp[4738]*kernel[0]+tmp[4739]*kernel[1]+tmp[4740]*kernel[2]+tmp[4838]*kernel[3]+tmp[4839]*kernel[4]+tmp[4840]*kernel[5]+tmp[4938]*kernel[6]+tmp[4939]*kernel[7]+tmp[4940]*kernel[8];
				ans[4840]<=tmp[4739]*kernel[0]+tmp[4740]*kernel[1]+tmp[4741]*kernel[2]+tmp[4839]*kernel[3]+tmp[4840]*kernel[4]+tmp[4841]*kernel[5]+tmp[4939]*kernel[6]+tmp[4940]*kernel[7]+tmp[4941]*kernel[8];
				ans[4841]<=tmp[4740]*kernel[0]+tmp[4741]*kernel[1]+tmp[4742]*kernel[2]+tmp[4840]*kernel[3]+tmp[4841]*kernel[4]+tmp[4842]*kernel[5]+tmp[4940]*kernel[6]+tmp[4941]*kernel[7]+tmp[4942]*kernel[8];
				ans[4842]<=tmp[4741]*kernel[0]+tmp[4742]*kernel[1]+tmp[4743]*kernel[2]+tmp[4841]*kernel[3]+tmp[4842]*kernel[4]+tmp[4843]*kernel[5]+tmp[4941]*kernel[6]+tmp[4942]*kernel[7]+tmp[4943]*kernel[8];
				ans[4843]<=tmp[4742]*kernel[0]+tmp[4743]*kernel[1]+tmp[4744]*kernel[2]+tmp[4842]*kernel[3]+tmp[4843]*kernel[4]+tmp[4844]*kernel[5]+tmp[4942]*kernel[6]+tmp[4943]*kernel[7]+tmp[4944]*kernel[8];
				ans[4844]<=tmp[4743]*kernel[0]+tmp[4744]*kernel[1]+tmp[4745]*kernel[2]+tmp[4843]*kernel[3]+tmp[4844]*kernel[4]+tmp[4845]*kernel[5]+tmp[4943]*kernel[6]+tmp[4944]*kernel[7]+tmp[4945]*kernel[8];
				ans[4845]<=tmp[4744]*kernel[0]+tmp[4745]*kernel[1]+tmp[4746]*kernel[2]+tmp[4844]*kernel[3]+tmp[4845]*kernel[4]+tmp[4846]*kernel[5]+tmp[4944]*kernel[6]+tmp[4945]*kernel[7]+tmp[4946]*kernel[8];
				ans[4846]<=tmp[4745]*kernel[0]+tmp[4746]*kernel[1]+tmp[4747]*kernel[2]+tmp[4845]*kernel[3]+tmp[4846]*kernel[4]+tmp[4847]*kernel[5]+tmp[4945]*kernel[6]+tmp[4946]*kernel[7]+tmp[4947]*kernel[8];
				ans[4847]<=tmp[4746]*kernel[0]+tmp[4747]*kernel[1]+tmp[4748]*kernel[2]+tmp[4846]*kernel[3]+tmp[4847]*kernel[4]+tmp[4848]*kernel[5]+tmp[4946]*kernel[6]+tmp[4947]*kernel[7]+tmp[4948]*kernel[8];
				ans[4848]<=tmp[4747]*kernel[0]+tmp[4748]*kernel[1]+tmp[4749]*kernel[2]+tmp[4847]*kernel[3]+tmp[4848]*kernel[4]+tmp[4849]*kernel[5]+tmp[4947]*kernel[6]+tmp[4948]*kernel[7]+tmp[4949]*kernel[8];
				ans[4849]<=tmp[4748]*kernel[0]+tmp[4749]*kernel[1]+tmp[4750]*kernel[2]+tmp[4848]*kernel[3]+tmp[4849]*kernel[4]+tmp[4850]*kernel[5]+tmp[4948]*kernel[6]+tmp[4949]*kernel[7]+tmp[4950]*kernel[8];
				ans[4850]<=tmp[4749]*kernel[0]+tmp[4750]*kernel[1]+tmp[4751]*kernel[2]+tmp[4849]*kernel[3]+tmp[4850]*kernel[4]+tmp[4851]*kernel[5]+tmp[4949]*kernel[6]+tmp[4950]*kernel[7]+tmp[4951]*kernel[8];
				ans[4851]<=tmp[4750]*kernel[0]+tmp[4751]*kernel[1]+tmp[4752]*kernel[2]+tmp[4850]*kernel[3]+tmp[4851]*kernel[4]+tmp[4852]*kernel[5]+tmp[4950]*kernel[6]+tmp[4951]*kernel[7]+tmp[4952]*kernel[8];
				ans[4852]<=tmp[4751]*kernel[0]+tmp[4752]*kernel[1]+tmp[4753]*kernel[2]+tmp[4851]*kernel[3]+tmp[4852]*kernel[4]+tmp[4853]*kernel[5]+tmp[4951]*kernel[6]+tmp[4952]*kernel[7]+tmp[4953]*kernel[8];
				ans[4853]<=tmp[4752]*kernel[0]+tmp[4753]*kernel[1]+tmp[4754]*kernel[2]+tmp[4852]*kernel[3]+tmp[4853]*kernel[4]+tmp[4854]*kernel[5]+tmp[4952]*kernel[6]+tmp[4953]*kernel[7]+tmp[4954]*kernel[8];
				ans[4854]<=tmp[4753]*kernel[0]+tmp[4754]*kernel[1]+tmp[4755]*kernel[2]+tmp[4853]*kernel[3]+tmp[4854]*kernel[4]+tmp[4855]*kernel[5]+tmp[4953]*kernel[6]+tmp[4954]*kernel[7]+tmp[4955]*kernel[8];
				ans[4855]<=tmp[4754]*kernel[0]+tmp[4755]*kernel[1]+tmp[4756]*kernel[2]+tmp[4854]*kernel[3]+tmp[4855]*kernel[4]+tmp[4856]*kernel[5]+tmp[4954]*kernel[6]+tmp[4955]*kernel[7]+tmp[4956]*kernel[8];
				ans[4856]<=tmp[4755]*kernel[0]+tmp[4756]*kernel[1]+tmp[4757]*kernel[2]+tmp[4855]*kernel[3]+tmp[4856]*kernel[4]+tmp[4857]*kernel[5]+tmp[4955]*kernel[6]+tmp[4956]*kernel[7]+tmp[4957]*kernel[8];
				ans[4857]<=tmp[4756]*kernel[0]+tmp[4757]*kernel[1]+tmp[4758]*kernel[2]+tmp[4856]*kernel[3]+tmp[4857]*kernel[4]+tmp[4858]*kernel[5]+tmp[4956]*kernel[6]+tmp[4957]*kernel[7]+tmp[4958]*kernel[8];
				ans[4858]<=tmp[4757]*kernel[0]+tmp[4758]*kernel[1]+tmp[4759]*kernel[2]+tmp[4857]*kernel[3]+tmp[4858]*kernel[4]+tmp[4859]*kernel[5]+tmp[4957]*kernel[6]+tmp[4958]*kernel[7]+tmp[4959]*kernel[8];
				ans[4859]<=tmp[4758]*kernel[0]+tmp[4759]*kernel[1]+tmp[4760]*kernel[2]+tmp[4858]*kernel[3]+tmp[4859]*kernel[4]+tmp[4860]*kernel[5]+tmp[4958]*kernel[6]+tmp[4959]*kernel[7]+tmp[4960]*kernel[8];
				ans[4860]<=tmp[4759]*kernel[0]+tmp[4760]*kernel[1]+tmp[4761]*kernel[2]+tmp[4859]*kernel[3]+tmp[4860]*kernel[4]+tmp[4861]*kernel[5]+tmp[4959]*kernel[6]+tmp[4960]*kernel[7]+tmp[4961]*kernel[8];
				ans[4861]<=tmp[4760]*kernel[0]+tmp[4761]*kernel[1]+tmp[4762]*kernel[2]+tmp[4860]*kernel[3]+tmp[4861]*kernel[4]+tmp[4862]*kernel[5]+tmp[4960]*kernel[6]+tmp[4961]*kernel[7]+tmp[4962]*kernel[8];
				ans[4862]<=tmp[4761]*kernel[0]+tmp[4762]*kernel[1]+tmp[4763]*kernel[2]+tmp[4861]*kernel[3]+tmp[4862]*kernel[4]+tmp[4863]*kernel[5]+tmp[4961]*kernel[6]+tmp[4962]*kernel[7]+tmp[4963]*kernel[8];
				ans[4863]<=tmp[4762]*kernel[0]+tmp[4763]*kernel[1]+tmp[4764]*kernel[2]+tmp[4862]*kernel[3]+tmp[4863]*kernel[4]+tmp[4864]*kernel[5]+tmp[4962]*kernel[6]+tmp[4963]*kernel[7]+tmp[4964]*kernel[8];
				ans[4864]<=tmp[4763]*kernel[0]+tmp[4764]*kernel[1]+tmp[4765]*kernel[2]+tmp[4863]*kernel[3]+tmp[4864]*kernel[4]+tmp[4865]*kernel[5]+tmp[4963]*kernel[6]+tmp[4964]*kernel[7]+tmp[4965]*kernel[8];
				ans[4865]<=tmp[4764]*kernel[0]+tmp[4765]*kernel[1]+tmp[4766]*kernel[2]+tmp[4864]*kernel[3]+tmp[4865]*kernel[4]+tmp[4866]*kernel[5]+tmp[4964]*kernel[6]+tmp[4965]*kernel[7]+tmp[4966]*kernel[8];
				ans[4866]<=tmp[4765]*kernel[0]+tmp[4766]*kernel[1]+tmp[4767]*kernel[2]+tmp[4865]*kernel[3]+tmp[4866]*kernel[4]+tmp[4867]*kernel[5]+tmp[4965]*kernel[6]+tmp[4966]*kernel[7]+tmp[4967]*kernel[8];
				ans[4867]<=tmp[4766]*kernel[0]+tmp[4767]*kernel[1]+tmp[4768]*kernel[2]+tmp[4866]*kernel[3]+tmp[4867]*kernel[4]+tmp[4868]*kernel[5]+tmp[4966]*kernel[6]+tmp[4967]*kernel[7]+tmp[4968]*kernel[8];
				ans[4868]<=tmp[4767]*kernel[0]+tmp[4768]*kernel[1]+tmp[4769]*kernel[2]+tmp[4867]*kernel[3]+tmp[4868]*kernel[4]+tmp[4869]*kernel[5]+tmp[4967]*kernel[6]+tmp[4968]*kernel[7]+tmp[4969]*kernel[8];
				ans[4869]<=tmp[4768]*kernel[0]+tmp[4769]*kernel[1]+tmp[4770]*kernel[2]+tmp[4868]*kernel[3]+tmp[4869]*kernel[4]+tmp[4870]*kernel[5]+tmp[4968]*kernel[6]+tmp[4969]*kernel[7]+tmp[4970]*kernel[8];
				ans[4870]<=tmp[4769]*kernel[0]+tmp[4770]*kernel[1]+tmp[4771]*kernel[2]+tmp[4869]*kernel[3]+tmp[4870]*kernel[4]+tmp[4871]*kernel[5]+tmp[4969]*kernel[6]+tmp[4970]*kernel[7]+tmp[4971]*kernel[8];
				ans[4871]<=tmp[4770]*kernel[0]+tmp[4771]*kernel[1]+tmp[4772]*kernel[2]+tmp[4870]*kernel[3]+tmp[4871]*kernel[4]+tmp[4872]*kernel[5]+tmp[4970]*kernel[6]+tmp[4971]*kernel[7]+tmp[4972]*kernel[8];
				ans[4872]<=tmp[4771]*kernel[0]+tmp[4772]*kernel[1]+tmp[4773]*kernel[2]+tmp[4871]*kernel[3]+tmp[4872]*kernel[4]+tmp[4873]*kernel[5]+tmp[4971]*kernel[6]+tmp[4972]*kernel[7]+tmp[4973]*kernel[8];
				ans[4873]<=tmp[4772]*kernel[0]+tmp[4773]*kernel[1]+tmp[4774]*kernel[2]+tmp[4872]*kernel[3]+tmp[4873]*kernel[4]+tmp[4874]*kernel[5]+tmp[4972]*kernel[6]+tmp[4973]*kernel[7]+tmp[4974]*kernel[8];
				ans[4874]<=tmp[4773]*kernel[0]+tmp[4774]*kernel[1]+tmp[4775]*kernel[2]+tmp[4873]*kernel[3]+tmp[4874]*kernel[4]+tmp[4875]*kernel[5]+tmp[4973]*kernel[6]+tmp[4974]*kernel[7]+tmp[4975]*kernel[8];
				ans[4875]<=tmp[4774]*kernel[0]+tmp[4775]*kernel[1]+tmp[4776]*kernel[2]+tmp[4874]*kernel[3]+tmp[4875]*kernel[4]+tmp[4876]*kernel[5]+tmp[4974]*kernel[6]+tmp[4975]*kernel[7]+tmp[4976]*kernel[8];
				ans[4876]<=tmp[4775]*kernel[0]+tmp[4776]*kernel[1]+tmp[4777]*kernel[2]+tmp[4875]*kernel[3]+tmp[4876]*kernel[4]+tmp[4877]*kernel[5]+tmp[4975]*kernel[6]+tmp[4976]*kernel[7]+tmp[4977]*kernel[8];
				ans[4877]<=tmp[4776]*kernel[0]+tmp[4777]*kernel[1]+tmp[4778]*kernel[2]+tmp[4876]*kernel[3]+tmp[4877]*kernel[4]+tmp[4878]*kernel[5]+tmp[4976]*kernel[6]+tmp[4977]*kernel[7]+tmp[4978]*kernel[8];
				ans[4878]<=tmp[4777]*kernel[0]+tmp[4778]*kernel[1]+tmp[4779]*kernel[2]+tmp[4877]*kernel[3]+tmp[4878]*kernel[4]+tmp[4879]*kernel[5]+tmp[4977]*kernel[6]+tmp[4978]*kernel[7]+tmp[4979]*kernel[8];
				ans[4879]<=tmp[4778]*kernel[0]+tmp[4779]*kernel[1]+tmp[4780]*kernel[2]+tmp[4878]*kernel[3]+tmp[4879]*kernel[4]+tmp[4880]*kernel[5]+tmp[4978]*kernel[6]+tmp[4979]*kernel[7]+tmp[4980]*kernel[8];
				ans[4880]<=tmp[4779]*kernel[0]+tmp[4780]*kernel[1]+tmp[4781]*kernel[2]+tmp[4879]*kernel[3]+tmp[4880]*kernel[4]+tmp[4881]*kernel[5]+tmp[4979]*kernel[6]+tmp[4980]*kernel[7]+tmp[4981]*kernel[8];
				ans[4881]<=tmp[4780]*kernel[0]+tmp[4781]*kernel[1]+tmp[4782]*kernel[2]+tmp[4880]*kernel[3]+tmp[4881]*kernel[4]+tmp[4882]*kernel[5]+tmp[4980]*kernel[6]+tmp[4981]*kernel[7]+tmp[4982]*kernel[8];
				ans[4882]<=tmp[4781]*kernel[0]+tmp[4782]*kernel[1]+tmp[4783]*kernel[2]+tmp[4881]*kernel[3]+tmp[4882]*kernel[4]+tmp[4883]*kernel[5]+tmp[4981]*kernel[6]+tmp[4982]*kernel[7]+tmp[4983]*kernel[8];
				ans[4883]<=tmp[4782]*kernel[0]+tmp[4783]*kernel[1]+tmp[4784]*kernel[2]+tmp[4882]*kernel[3]+tmp[4883]*kernel[4]+tmp[4884]*kernel[5]+tmp[4982]*kernel[6]+tmp[4983]*kernel[7]+tmp[4984]*kernel[8];
				ans[4884]<=tmp[4783]*kernel[0]+tmp[4784]*kernel[1]+tmp[4785]*kernel[2]+tmp[4883]*kernel[3]+tmp[4884]*kernel[4]+tmp[4885]*kernel[5]+tmp[4983]*kernel[6]+tmp[4984]*kernel[7]+tmp[4985]*kernel[8];
				ans[4885]<=tmp[4784]*kernel[0]+tmp[4785]*kernel[1]+tmp[4786]*kernel[2]+tmp[4884]*kernel[3]+tmp[4885]*kernel[4]+tmp[4886]*kernel[5]+tmp[4984]*kernel[6]+tmp[4985]*kernel[7]+tmp[4986]*kernel[8];
				ans[4886]<=tmp[4785]*kernel[0]+tmp[4786]*kernel[1]+tmp[4787]*kernel[2]+tmp[4885]*kernel[3]+tmp[4886]*kernel[4]+tmp[4887]*kernel[5]+tmp[4985]*kernel[6]+tmp[4986]*kernel[7]+tmp[4987]*kernel[8];
				ans[4887]<=tmp[4786]*kernel[0]+tmp[4787]*kernel[1]+tmp[4788]*kernel[2]+tmp[4886]*kernel[3]+tmp[4887]*kernel[4]+tmp[4888]*kernel[5]+tmp[4986]*kernel[6]+tmp[4987]*kernel[7]+tmp[4988]*kernel[8];
				ans[4888]<=tmp[4787]*kernel[0]+tmp[4788]*kernel[1]+tmp[4789]*kernel[2]+tmp[4887]*kernel[3]+tmp[4888]*kernel[4]+tmp[4889]*kernel[5]+tmp[4987]*kernel[6]+tmp[4988]*kernel[7]+tmp[4989]*kernel[8];
				ans[4889]<=tmp[4788]*kernel[0]+tmp[4789]*kernel[1]+tmp[4790]*kernel[2]+tmp[4888]*kernel[3]+tmp[4889]*kernel[4]+tmp[4890]*kernel[5]+tmp[4988]*kernel[6]+tmp[4989]*kernel[7]+tmp[4990]*kernel[8];
				ans[4890]<=tmp[4789]*kernel[0]+tmp[4790]*kernel[1]+tmp[4791]*kernel[2]+tmp[4889]*kernel[3]+tmp[4890]*kernel[4]+tmp[4891]*kernel[5]+tmp[4989]*kernel[6]+tmp[4990]*kernel[7]+tmp[4991]*kernel[8];
				ans[4891]<=tmp[4790]*kernel[0]+tmp[4791]*kernel[1]+tmp[4792]*kernel[2]+tmp[4890]*kernel[3]+tmp[4891]*kernel[4]+tmp[4892]*kernel[5]+tmp[4990]*kernel[6]+tmp[4991]*kernel[7]+tmp[4992]*kernel[8];
				ans[4892]<=tmp[4791]*kernel[0]+tmp[4792]*kernel[1]+tmp[4793]*kernel[2]+tmp[4891]*kernel[3]+tmp[4892]*kernel[4]+tmp[4893]*kernel[5]+tmp[4991]*kernel[6]+tmp[4992]*kernel[7]+tmp[4993]*kernel[8];
				ans[4893]<=tmp[4792]*kernel[0]+tmp[4793]*kernel[1]+tmp[4794]*kernel[2]+tmp[4892]*kernel[3]+tmp[4893]*kernel[4]+tmp[4894]*kernel[5]+tmp[4992]*kernel[6]+tmp[4993]*kernel[7]+tmp[4994]*kernel[8];
				ans[4894]<=tmp[4793]*kernel[0]+tmp[4794]*kernel[1]+tmp[4795]*kernel[2]+tmp[4893]*kernel[3]+tmp[4894]*kernel[4]+tmp[4895]*kernel[5]+tmp[4993]*kernel[6]+tmp[4994]*kernel[7]+tmp[4995]*kernel[8];
				ans[4895]<=tmp[4794]*kernel[0]+tmp[4795]*kernel[1]+tmp[4796]*kernel[2]+tmp[4894]*kernel[3]+tmp[4895]*kernel[4]+tmp[4896]*kernel[5]+tmp[4994]*kernel[6]+tmp[4995]*kernel[7]+tmp[4996]*kernel[8];
				ans[4896]<=tmp[4795]*kernel[0]+tmp[4796]*kernel[1]+tmp[4797]*kernel[2]+tmp[4895]*kernel[3]+tmp[4896]*kernel[4]+tmp[4897]*kernel[5]+tmp[4995]*kernel[6]+tmp[4996]*kernel[7]+tmp[4997]*kernel[8];
				ans[4897]<=tmp[4796]*kernel[0]+tmp[4797]*kernel[1]+tmp[4798]*kernel[2]+tmp[4896]*kernel[3]+tmp[4897]*kernel[4]+tmp[4898]*kernel[5]+tmp[4996]*kernel[6]+tmp[4997]*kernel[7]+tmp[4998]*kernel[8];
				ans[4898]<=tmp[4797]*kernel[0]+tmp[4798]*kernel[1]+tmp[4799]*kernel[2]+tmp[4897]*kernel[3]+tmp[4898]*kernel[4]+tmp[4899]*kernel[5]+tmp[4997]*kernel[6]+tmp[4998]*kernel[7]+tmp[4999]*kernel[8];
				ans[4899]<=tmp[4798]*kernel[0]+tmp[4799]*kernel[1]+tmp[4898]*kernel[3]+tmp[4899]*kernel[4]+tmp[4998]*kernel[6]+tmp[4999]*kernel[7];
				ans[4900]<=tmp[4800]*kernel[1]+tmp[4801]*kernel[2]+tmp[4900]*kernel[4]+tmp[4901]*kernel[5]+tmp[5000]*kernel[7]+tmp[5001]*kernel[8];
				ans[4901]<=tmp[4800]*kernel[0]+tmp[4801]*kernel[1]+tmp[4802]*kernel[2]+tmp[4900]*kernel[3]+tmp[4901]*kernel[4]+tmp[4902]*kernel[5]+tmp[5000]*kernel[6]+tmp[5001]*kernel[7]+tmp[5002]*kernel[8];
				ans[4902]<=tmp[4801]*kernel[0]+tmp[4802]*kernel[1]+tmp[4803]*kernel[2]+tmp[4901]*kernel[3]+tmp[4902]*kernel[4]+tmp[4903]*kernel[5]+tmp[5001]*kernel[6]+tmp[5002]*kernel[7]+tmp[5003]*kernel[8];
				ans[4903]<=tmp[4802]*kernel[0]+tmp[4803]*kernel[1]+tmp[4804]*kernel[2]+tmp[4902]*kernel[3]+tmp[4903]*kernel[4]+tmp[4904]*kernel[5]+tmp[5002]*kernel[6]+tmp[5003]*kernel[7]+tmp[5004]*kernel[8];
				ans[4904]<=tmp[4803]*kernel[0]+tmp[4804]*kernel[1]+tmp[4805]*kernel[2]+tmp[4903]*kernel[3]+tmp[4904]*kernel[4]+tmp[4905]*kernel[5]+tmp[5003]*kernel[6]+tmp[5004]*kernel[7]+tmp[5005]*kernel[8];
				ans[4905]<=tmp[4804]*kernel[0]+tmp[4805]*kernel[1]+tmp[4806]*kernel[2]+tmp[4904]*kernel[3]+tmp[4905]*kernel[4]+tmp[4906]*kernel[5]+tmp[5004]*kernel[6]+tmp[5005]*kernel[7]+tmp[5006]*kernel[8];
				ans[4906]<=tmp[4805]*kernel[0]+tmp[4806]*kernel[1]+tmp[4807]*kernel[2]+tmp[4905]*kernel[3]+tmp[4906]*kernel[4]+tmp[4907]*kernel[5]+tmp[5005]*kernel[6]+tmp[5006]*kernel[7]+tmp[5007]*kernel[8];
				ans[4907]<=tmp[4806]*kernel[0]+tmp[4807]*kernel[1]+tmp[4808]*kernel[2]+tmp[4906]*kernel[3]+tmp[4907]*kernel[4]+tmp[4908]*kernel[5]+tmp[5006]*kernel[6]+tmp[5007]*kernel[7]+tmp[5008]*kernel[8];
				ans[4908]<=tmp[4807]*kernel[0]+tmp[4808]*kernel[1]+tmp[4809]*kernel[2]+tmp[4907]*kernel[3]+tmp[4908]*kernel[4]+tmp[4909]*kernel[5]+tmp[5007]*kernel[6]+tmp[5008]*kernel[7]+tmp[5009]*kernel[8];
				ans[4909]<=tmp[4808]*kernel[0]+tmp[4809]*kernel[1]+tmp[4810]*kernel[2]+tmp[4908]*kernel[3]+tmp[4909]*kernel[4]+tmp[4910]*kernel[5]+tmp[5008]*kernel[6]+tmp[5009]*kernel[7]+tmp[5010]*kernel[8];
				ans[4910]<=tmp[4809]*kernel[0]+tmp[4810]*kernel[1]+tmp[4811]*kernel[2]+tmp[4909]*kernel[3]+tmp[4910]*kernel[4]+tmp[4911]*kernel[5]+tmp[5009]*kernel[6]+tmp[5010]*kernel[7]+tmp[5011]*kernel[8];
				ans[4911]<=tmp[4810]*kernel[0]+tmp[4811]*kernel[1]+tmp[4812]*kernel[2]+tmp[4910]*kernel[3]+tmp[4911]*kernel[4]+tmp[4912]*kernel[5]+tmp[5010]*kernel[6]+tmp[5011]*kernel[7]+tmp[5012]*kernel[8];
				ans[4912]<=tmp[4811]*kernel[0]+tmp[4812]*kernel[1]+tmp[4813]*kernel[2]+tmp[4911]*kernel[3]+tmp[4912]*kernel[4]+tmp[4913]*kernel[5]+tmp[5011]*kernel[6]+tmp[5012]*kernel[7]+tmp[5013]*kernel[8];
				ans[4913]<=tmp[4812]*kernel[0]+tmp[4813]*kernel[1]+tmp[4814]*kernel[2]+tmp[4912]*kernel[3]+tmp[4913]*kernel[4]+tmp[4914]*kernel[5]+tmp[5012]*kernel[6]+tmp[5013]*kernel[7]+tmp[5014]*kernel[8];
				ans[4914]<=tmp[4813]*kernel[0]+tmp[4814]*kernel[1]+tmp[4815]*kernel[2]+tmp[4913]*kernel[3]+tmp[4914]*kernel[4]+tmp[4915]*kernel[5]+tmp[5013]*kernel[6]+tmp[5014]*kernel[7]+tmp[5015]*kernel[8];
				ans[4915]<=tmp[4814]*kernel[0]+tmp[4815]*kernel[1]+tmp[4816]*kernel[2]+tmp[4914]*kernel[3]+tmp[4915]*kernel[4]+tmp[4916]*kernel[5]+tmp[5014]*kernel[6]+tmp[5015]*kernel[7]+tmp[5016]*kernel[8];
				ans[4916]<=tmp[4815]*kernel[0]+tmp[4816]*kernel[1]+tmp[4817]*kernel[2]+tmp[4915]*kernel[3]+tmp[4916]*kernel[4]+tmp[4917]*kernel[5]+tmp[5015]*kernel[6]+tmp[5016]*kernel[7]+tmp[5017]*kernel[8];
				ans[4917]<=tmp[4816]*kernel[0]+tmp[4817]*kernel[1]+tmp[4818]*kernel[2]+tmp[4916]*kernel[3]+tmp[4917]*kernel[4]+tmp[4918]*kernel[5]+tmp[5016]*kernel[6]+tmp[5017]*kernel[7]+tmp[5018]*kernel[8];
				ans[4918]<=tmp[4817]*kernel[0]+tmp[4818]*kernel[1]+tmp[4819]*kernel[2]+tmp[4917]*kernel[3]+tmp[4918]*kernel[4]+tmp[4919]*kernel[5]+tmp[5017]*kernel[6]+tmp[5018]*kernel[7]+tmp[5019]*kernel[8];
				ans[4919]<=tmp[4818]*kernel[0]+tmp[4819]*kernel[1]+tmp[4820]*kernel[2]+tmp[4918]*kernel[3]+tmp[4919]*kernel[4]+tmp[4920]*kernel[5]+tmp[5018]*kernel[6]+tmp[5019]*kernel[7]+tmp[5020]*kernel[8];
				ans[4920]<=tmp[4819]*kernel[0]+tmp[4820]*kernel[1]+tmp[4821]*kernel[2]+tmp[4919]*kernel[3]+tmp[4920]*kernel[4]+tmp[4921]*kernel[5]+tmp[5019]*kernel[6]+tmp[5020]*kernel[7]+tmp[5021]*kernel[8];
				ans[4921]<=tmp[4820]*kernel[0]+tmp[4821]*kernel[1]+tmp[4822]*kernel[2]+tmp[4920]*kernel[3]+tmp[4921]*kernel[4]+tmp[4922]*kernel[5]+tmp[5020]*kernel[6]+tmp[5021]*kernel[7]+tmp[5022]*kernel[8];
				ans[4922]<=tmp[4821]*kernel[0]+tmp[4822]*kernel[1]+tmp[4823]*kernel[2]+tmp[4921]*kernel[3]+tmp[4922]*kernel[4]+tmp[4923]*kernel[5]+tmp[5021]*kernel[6]+tmp[5022]*kernel[7]+tmp[5023]*kernel[8];
				ans[4923]<=tmp[4822]*kernel[0]+tmp[4823]*kernel[1]+tmp[4824]*kernel[2]+tmp[4922]*kernel[3]+tmp[4923]*kernel[4]+tmp[4924]*kernel[5]+tmp[5022]*kernel[6]+tmp[5023]*kernel[7]+tmp[5024]*kernel[8];
				ans[4924]<=tmp[4823]*kernel[0]+tmp[4824]*kernel[1]+tmp[4825]*kernel[2]+tmp[4923]*kernel[3]+tmp[4924]*kernel[4]+tmp[4925]*kernel[5]+tmp[5023]*kernel[6]+tmp[5024]*kernel[7]+tmp[5025]*kernel[8];
				ans[4925]<=tmp[4824]*kernel[0]+tmp[4825]*kernel[1]+tmp[4826]*kernel[2]+tmp[4924]*kernel[3]+tmp[4925]*kernel[4]+tmp[4926]*kernel[5]+tmp[5024]*kernel[6]+tmp[5025]*kernel[7]+tmp[5026]*kernel[8];
				ans[4926]<=tmp[4825]*kernel[0]+tmp[4826]*kernel[1]+tmp[4827]*kernel[2]+tmp[4925]*kernel[3]+tmp[4926]*kernel[4]+tmp[4927]*kernel[5]+tmp[5025]*kernel[6]+tmp[5026]*kernel[7]+tmp[5027]*kernel[8];
				ans[4927]<=tmp[4826]*kernel[0]+tmp[4827]*kernel[1]+tmp[4828]*kernel[2]+tmp[4926]*kernel[3]+tmp[4927]*kernel[4]+tmp[4928]*kernel[5]+tmp[5026]*kernel[6]+tmp[5027]*kernel[7]+tmp[5028]*kernel[8];
				ans[4928]<=tmp[4827]*kernel[0]+tmp[4828]*kernel[1]+tmp[4829]*kernel[2]+tmp[4927]*kernel[3]+tmp[4928]*kernel[4]+tmp[4929]*kernel[5]+tmp[5027]*kernel[6]+tmp[5028]*kernel[7]+tmp[5029]*kernel[8];
				ans[4929]<=tmp[4828]*kernel[0]+tmp[4829]*kernel[1]+tmp[4830]*kernel[2]+tmp[4928]*kernel[3]+tmp[4929]*kernel[4]+tmp[4930]*kernel[5]+tmp[5028]*kernel[6]+tmp[5029]*kernel[7]+tmp[5030]*kernel[8];
				ans[4930]<=tmp[4829]*kernel[0]+tmp[4830]*kernel[1]+tmp[4831]*kernel[2]+tmp[4929]*kernel[3]+tmp[4930]*kernel[4]+tmp[4931]*kernel[5]+tmp[5029]*kernel[6]+tmp[5030]*kernel[7]+tmp[5031]*kernel[8];
				ans[4931]<=tmp[4830]*kernel[0]+tmp[4831]*kernel[1]+tmp[4832]*kernel[2]+tmp[4930]*kernel[3]+tmp[4931]*kernel[4]+tmp[4932]*kernel[5]+tmp[5030]*kernel[6]+tmp[5031]*kernel[7]+tmp[5032]*kernel[8];
				ans[4932]<=tmp[4831]*kernel[0]+tmp[4832]*kernel[1]+tmp[4833]*kernel[2]+tmp[4931]*kernel[3]+tmp[4932]*kernel[4]+tmp[4933]*kernel[5]+tmp[5031]*kernel[6]+tmp[5032]*kernel[7]+tmp[5033]*kernel[8];
				ans[4933]<=tmp[4832]*kernel[0]+tmp[4833]*kernel[1]+tmp[4834]*kernel[2]+tmp[4932]*kernel[3]+tmp[4933]*kernel[4]+tmp[4934]*kernel[5]+tmp[5032]*kernel[6]+tmp[5033]*kernel[7]+tmp[5034]*kernel[8];
				ans[4934]<=tmp[4833]*kernel[0]+tmp[4834]*kernel[1]+tmp[4835]*kernel[2]+tmp[4933]*kernel[3]+tmp[4934]*kernel[4]+tmp[4935]*kernel[5]+tmp[5033]*kernel[6]+tmp[5034]*kernel[7]+tmp[5035]*kernel[8];
				ans[4935]<=tmp[4834]*kernel[0]+tmp[4835]*kernel[1]+tmp[4836]*kernel[2]+tmp[4934]*kernel[3]+tmp[4935]*kernel[4]+tmp[4936]*kernel[5]+tmp[5034]*kernel[6]+tmp[5035]*kernel[7]+tmp[5036]*kernel[8];
				ans[4936]<=tmp[4835]*kernel[0]+tmp[4836]*kernel[1]+tmp[4837]*kernel[2]+tmp[4935]*kernel[3]+tmp[4936]*kernel[4]+tmp[4937]*kernel[5]+tmp[5035]*kernel[6]+tmp[5036]*kernel[7]+tmp[5037]*kernel[8];
				ans[4937]<=tmp[4836]*kernel[0]+tmp[4837]*kernel[1]+tmp[4838]*kernel[2]+tmp[4936]*kernel[3]+tmp[4937]*kernel[4]+tmp[4938]*kernel[5]+tmp[5036]*kernel[6]+tmp[5037]*kernel[7]+tmp[5038]*kernel[8];
				ans[4938]<=tmp[4837]*kernel[0]+tmp[4838]*kernel[1]+tmp[4839]*kernel[2]+tmp[4937]*kernel[3]+tmp[4938]*kernel[4]+tmp[4939]*kernel[5]+tmp[5037]*kernel[6]+tmp[5038]*kernel[7]+tmp[5039]*kernel[8];
				ans[4939]<=tmp[4838]*kernel[0]+tmp[4839]*kernel[1]+tmp[4840]*kernel[2]+tmp[4938]*kernel[3]+tmp[4939]*kernel[4]+tmp[4940]*kernel[5]+tmp[5038]*kernel[6]+tmp[5039]*kernel[7]+tmp[5040]*kernel[8];
				ans[4940]<=tmp[4839]*kernel[0]+tmp[4840]*kernel[1]+tmp[4841]*kernel[2]+tmp[4939]*kernel[3]+tmp[4940]*kernel[4]+tmp[4941]*kernel[5]+tmp[5039]*kernel[6]+tmp[5040]*kernel[7]+tmp[5041]*kernel[8];
				ans[4941]<=tmp[4840]*kernel[0]+tmp[4841]*kernel[1]+tmp[4842]*kernel[2]+tmp[4940]*kernel[3]+tmp[4941]*kernel[4]+tmp[4942]*kernel[5]+tmp[5040]*kernel[6]+tmp[5041]*kernel[7]+tmp[5042]*kernel[8];
				ans[4942]<=tmp[4841]*kernel[0]+tmp[4842]*kernel[1]+tmp[4843]*kernel[2]+tmp[4941]*kernel[3]+tmp[4942]*kernel[4]+tmp[4943]*kernel[5]+tmp[5041]*kernel[6]+tmp[5042]*kernel[7]+tmp[5043]*kernel[8];
				ans[4943]<=tmp[4842]*kernel[0]+tmp[4843]*kernel[1]+tmp[4844]*kernel[2]+tmp[4942]*kernel[3]+tmp[4943]*kernel[4]+tmp[4944]*kernel[5]+tmp[5042]*kernel[6]+tmp[5043]*kernel[7]+tmp[5044]*kernel[8];
				ans[4944]<=tmp[4843]*kernel[0]+tmp[4844]*kernel[1]+tmp[4845]*kernel[2]+tmp[4943]*kernel[3]+tmp[4944]*kernel[4]+tmp[4945]*kernel[5]+tmp[5043]*kernel[6]+tmp[5044]*kernel[7]+tmp[5045]*kernel[8];
				ans[4945]<=tmp[4844]*kernel[0]+tmp[4845]*kernel[1]+tmp[4846]*kernel[2]+tmp[4944]*kernel[3]+tmp[4945]*kernel[4]+tmp[4946]*kernel[5]+tmp[5044]*kernel[6]+tmp[5045]*kernel[7]+tmp[5046]*kernel[8];
				ans[4946]<=tmp[4845]*kernel[0]+tmp[4846]*kernel[1]+tmp[4847]*kernel[2]+tmp[4945]*kernel[3]+tmp[4946]*kernel[4]+tmp[4947]*kernel[5]+tmp[5045]*kernel[6]+tmp[5046]*kernel[7]+tmp[5047]*kernel[8];
				ans[4947]<=tmp[4846]*kernel[0]+tmp[4847]*kernel[1]+tmp[4848]*kernel[2]+tmp[4946]*kernel[3]+tmp[4947]*kernel[4]+tmp[4948]*kernel[5]+tmp[5046]*kernel[6]+tmp[5047]*kernel[7]+tmp[5048]*kernel[8];
				ans[4948]<=tmp[4847]*kernel[0]+tmp[4848]*kernel[1]+tmp[4849]*kernel[2]+tmp[4947]*kernel[3]+tmp[4948]*kernel[4]+tmp[4949]*kernel[5]+tmp[5047]*kernel[6]+tmp[5048]*kernel[7]+tmp[5049]*kernel[8];
				ans[4949]<=tmp[4848]*kernel[0]+tmp[4849]*kernel[1]+tmp[4850]*kernel[2]+tmp[4948]*kernel[3]+tmp[4949]*kernel[4]+tmp[4950]*kernel[5]+tmp[5048]*kernel[6]+tmp[5049]*kernel[7]+tmp[5050]*kernel[8];
				ans[4950]<=tmp[4849]*kernel[0]+tmp[4850]*kernel[1]+tmp[4851]*kernel[2]+tmp[4949]*kernel[3]+tmp[4950]*kernel[4]+tmp[4951]*kernel[5]+tmp[5049]*kernel[6]+tmp[5050]*kernel[7]+tmp[5051]*kernel[8];
				ans[4951]<=tmp[4850]*kernel[0]+tmp[4851]*kernel[1]+tmp[4852]*kernel[2]+tmp[4950]*kernel[3]+tmp[4951]*kernel[4]+tmp[4952]*kernel[5]+tmp[5050]*kernel[6]+tmp[5051]*kernel[7]+tmp[5052]*kernel[8];
				ans[4952]<=tmp[4851]*kernel[0]+tmp[4852]*kernel[1]+tmp[4853]*kernel[2]+tmp[4951]*kernel[3]+tmp[4952]*kernel[4]+tmp[4953]*kernel[5]+tmp[5051]*kernel[6]+tmp[5052]*kernel[7]+tmp[5053]*kernel[8];
				ans[4953]<=tmp[4852]*kernel[0]+tmp[4853]*kernel[1]+tmp[4854]*kernel[2]+tmp[4952]*kernel[3]+tmp[4953]*kernel[4]+tmp[4954]*kernel[5]+tmp[5052]*kernel[6]+tmp[5053]*kernel[7]+tmp[5054]*kernel[8];
				ans[4954]<=tmp[4853]*kernel[0]+tmp[4854]*kernel[1]+tmp[4855]*kernel[2]+tmp[4953]*kernel[3]+tmp[4954]*kernel[4]+tmp[4955]*kernel[5]+tmp[5053]*kernel[6]+tmp[5054]*kernel[7]+tmp[5055]*kernel[8];
				ans[4955]<=tmp[4854]*kernel[0]+tmp[4855]*kernel[1]+tmp[4856]*kernel[2]+tmp[4954]*kernel[3]+tmp[4955]*kernel[4]+tmp[4956]*kernel[5]+tmp[5054]*kernel[6]+tmp[5055]*kernel[7]+tmp[5056]*kernel[8];
				ans[4956]<=tmp[4855]*kernel[0]+tmp[4856]*kernel[1]+tmp[4857]*kernel[2]+tmp[4955]*kernel[3]+tmp[4956]*kernel[4]+tmp[4957]*kernel[5]+tmp[5055]*kernel[6]+tmp[5056]*kernel[7]+tmp[5057]*kernel[8];
				ans[4957]<=tmp[4856]*kernel[0]+tmp[4857]*kernel[1]+tmp[4858]*kernel[2]+tmp[4956]*kernel[3]+tmp[4957]*kernel[4]+tmp[4958]*kernel[5]+tmp[5056]*kernel[6]+tmp[5057]*kernel[7]+tmp[5058]*kernel[8];
				ans[4958]<=tmp[4857]*kernel[0]+tmp[4858]*kernel[1]+tmp[4859]*kernel[2]+tmp[4957]*kernel[3]+tmp[4958]*kernel[4]+tmp[4959]*kernel[5]+tmp[5057]*kernel[6]+tmp[5058]*kernel[7]+tmp[5059]*kernel[8];
				ans[4959]<=tmp[4858]*kernel[0]+tmp[4859]*kernel[1]+tmp[4860]*kernel[2]+tmp[4958]*kernel[3]+tmp[4959]*kernel[4]+tmp[4960]*kernel[5]+tmp[5058]*kernel[6]+tmp[5059]*kernel[7]+tmp[5060]*kernel[8];
				ans[4960]<=tmp[4859]*kernel[0]+tmp[4860]*kernel[1]+tmp[4861]*kernel[2]+tmp[4959]*kernel[3]+tmp[4960]*kernel[4]+tmp[4961]*kernel[5]+tmp[5059]*kernel[6]+tmp[5060]*kernel[7]+tmp[5061]*kernel[8];
				ans[4961]<=tmp[4860]*kernel[0]+tmp[4861]*kernel[1]+tmp[4862]*kernel[2]+tmp[4960]*kernel[3]+tmp[4961]*kernel[4]+tmp[4962]*kernel[5]+tmp[5060]*kernel[6]+tmp[5061]*kernel[7]+tmp[5062]*kernel[8];
				ans[4962]<=tmp[4861]*kernel[0]+tmp[4862]*kernel[1]+tmp[4863]*kernel[2]+tmp[4961]*kernel[3]+tmp[4962]*kernel[4]+tmp[4963]*kernel[5]+tmp[5061]*kernel[6]+tmp[5062]*kernel[7]+tmp[5063]*kernel[8];
				ans[4963]<=tmp[4862]*kernel[0]+tmp[4863]*kernel[1]+tmp[4864]*kernel[2]+tmp[4962]*kernel[3]+tmp[4963]*kernel[4]+tmp[4964]*kernel[5]+tmp[5062]*kernel[6]+tmp[5063]*kernel[7]+tmp[5064]*kernel[8];
				ans[4964]<=tmp[4863]*kernel[0]+tmp[4864]*kernel[1]+tmp[4865]*kernel[2]+tmp[4963]*kernel[3]+tmp[4964]*kernel[4]+tmp[4965]*kernel[5]+tmp[5063]*kernel[6]+tmp[5064]*kernel[7]+tmp[5065]*kernel[8];
				ans[4965]<=tmp[4864]*kernel[0]+tmp[4865]*kernel[1]+tmp[4866]*kernel[2]+tmp[4964]*kernel[3]+tmp[4965]*kernel[4]+tmp[4966]*kernel[5]+tmp[5064]*kernel[6]+tmp[5065]*kernel[7]+tmp[5066]*kernel[8];
				ans[4966]<=tmp[4865]*kernel[0]+tmp[4866]*kernel[1]+tmp[4867]*kernel[2]+tmp[4965]*kernel[3]+tmp[4966]*kernel[4]+tmp[4967]*kernel[5]+tmp[5065]*kernel[6]+tmp[5066]*kernel[7]+tmp[5067]*kernel[8];
				ans[4967]<=tmp[4866]*kernel[0]+tmp[4867]*kernel[1]+tmp[4868]*kernel[2]+tmp[4966]*kernel[3]+tmp[4967]*kernel[4]+tmp[4968]*kernel[5]+tmp[5066]*kernel[6]+tmp[5067]*kernel[7]+tmp[5068]*kernel[8];
				ans[4968]<=tmp[4867]*kernel[0]+tmp[4868]*kernel[1]+tmp[4869]*kernel[2]+tmp[4967]*kernel[3]+tmp[4968]*kernel[4]+tmp[4969]*kernel[5]+tmp[5067]*kernel[6]+tmp[5068]*kernel[7]+tmp[5069]*kernel[8];
				ans[4969]<=tmp[4868]*kernel[0]+tmp[4869]*kernel[1]+tmp[4870]*kernel[2]+tmp[4968]*kernel[3]+tmp[4969]*kernel[4]+tmp[4970]*kernel[5]+tmp[5068]*kernel[6]+tmp[5069]*kernel[7]+tmp[5070]*kernel[8];
				ans[4970]<=tmp[4869]*kernel[0]+tmp[4870]*kernel[1]+tmp[4871]*kernel[2]+tmp[4969]*kernel[3]+tmp[4970]*kernel[4]+tmp[4971]*kernel[5]+tmp[5069]*kernel[6]+tmp[5070]*kernel[7]+tmp[5071]*kernel[8];
				ans[4971]<=tmp[4870]*kernel[0]+tmp[4871]*kernel[1]+tmp[4872]*kernel[2]+tmp[4970]*kernel[3]+tmp[4971]*kernel[4]+tmp[4972]*kernel[5]+tmp[5070]*kernel[6]+tmp[5071]*kernel[7]+tmp[5072]*kernel[8];
				ans[4972]<=tmp[4871]*kernel[0]+tmp[4872]*kernel[1]+tmp[4873]*kernel[2]+tmp[4971]*kernel[3]+tmp[4972]*kernel[4]+tmp[4973]*kernel[5]+tmp[5071]*kernel[6]+tmp[5072]*kernel[7]+tmp[5073]*kernel[8];
				ans[4973]<=tmp[4872]*kernel[0]+tmp[4873]*kernel[1]+tmp[4874]*kernel[2]+tmp[4972]*kernel[3]+tmp[4973]*kernel[4]+tmp[4974]*kernel[5]+tmp[5072]*kernel[6]+tmp[5073]*kernel[7]+tmp[5074]*kernel[8];
				ans[4974]<=tmp[4873]*kernel[0]+tmp[4874]*kernel[1]+tmp[4875]*kernel[2]+tmp[4973]*kernel[3]+tmp[4974]*kernel[4]+tmp[4975]*kernel[5]+tmp[5073]*kernel[6]+tmp[5074]*kernel[7]+tmp[5075]*kernel[8];
				ans[4975]<=tmp[4874]*kernel[0]+tmp[4875]*kernel[1]+tmp[4876]*kernel[2]+tmp[4974]*kernel[3]+tmp[4975]*kernel[4]+tmp[4976]*kernel[5]+tmp[5074]*kernel[6]+tmp[5075]*kernel[7]+tmp[5076]*kernel[8];
				ans[4976]<=tmp[4875]*kernel[0]+tmp[4876]*kernel[1]+tmp[4877]*kernel[2]+tmp[4975]*kernel[3]+tmp[4976]*kernel[4]+tmp[4977]*kernel[5]+tmp[5075]*kernel[6]+tmp[5076]*kernel[7]+tmp[5077]*kernel[8];
				ans[4977]<=tmp[4876]*kernel[0]+tmp[4877]*kernel[1]+tmp[4878]*kernel[2]+tmp[4976]*kernel[3]+tmp[4977]*kernel[4]+tmp[4978]*kernel[5]+tmp[5076]*kernel[6]+tmp[5077]*kernel[7]+tmp[5078]*kernel[8];
				ans[4978]<=tmp[4877]*kernel[0]+tmp[4878]*kernel[1]+tmp[4879]*kernel[2]+tmp[4977]*kernel[3]+tmp[4978]*kernel[4]+tmp[4979]*kernel[5]+tmp[5077]*kernel[6]+tmp[5078]*kernel[7]+tmp[5079]*kernel[8];
				ans[4979]<=tmp[4878]*kernel[0]+tmp[4879]*kernel[1]+tmp[4880]*kernel[2]+tmp[4978]*kernel[3]+tmp[4979]*kernel[4]+tmp[4980]*kernel[5]+tmp[5078]*kernel[6]+tmp[5079]*kernel[7]+tmp[5080]*kernel[8];
				ans[4980]<=tmp[4879]*kernel[0]+tmp[4880]*kernel[1]+tmp[4881]*kernel[2]+tmp[4979]*kernel[3]+tmp[4980]*kernel[4]+tmp[4981]*kernel[5]+tmp[5079]*kernel[6]+tmp[5080]*kernel[7]+tmp[5081]*kernel[8];
				ans[4981]<=tmp[4880]*kernel[0]+tmp[4881]*kernel[1]+tmp[4882]*kernel[2]+tmp[4980]*kernel[3]+tmp[4981]*kernel[4]+tmp[4982]*kernel[5]+tmp[5080]*kernel[6]+tmp[5081]*kernel[7]+tmp[5082]*kernel[8];
				ans[4982]<=tmp[4881]*kernel[0]+tmp[4882]*kernel[1]+tmp[4883]*kernel[2]+tmp[4981]*kernel[3]+tmp[4982]*kernel[4]+tmp[4983]*kernel[5]+tmp[5081]*kernel[6]+tmp[5082]*kernel[7]+tmp[5083]*kernel[8];
				ans[4983]<=tmp[4882]*kernel[0]+tmp[4883]*kernel[1]+tmp[4884]*kernel[2]+tmp[4982]*kernel[3]+tmp[4983]*kernel[4]+tmp[4984]*kernel[5]+tmp[5082]*kernel[6]+tmp[5083]*kernel[7]+tmp[5084]*kernel[8];
				ans[4984]<=tmp[4883]*kernel[0]+tmp[4884]*kernel[1]+tmp[4885]*kernel[2]+tmp[4983]*kernel[3]+tmp[4984]*kernel[4]+tmp[4985]*kernel[5]+tmp[5083]*kernel[6]+tmp[5084]*kernel[7]+tmp[5085]*kernel[8];
				ans[4985]<=tmp[4884]*kernel[0]+tmp[4885]*kernel[1]+tmp[4886]*kernel[2]+tmp[4984]*kernel[3]+tmp[4985]*kernel[4]+tmp[4986]*kernel[5]+tmp[5084]*kernel[6]+tmp[5085]*kernel[7]+tmp[5086]*kernel[8];
				ans[4986]<=tmp[4885]*kernel[0]+tmp[4886]*kernel[1]+tmp[4887]*kernel[2]+tmp[4985]*kernel[3]+tmp[4986]*kernel[4]+tmp[4987]*kernel[5]+tmp[5085]*kernel[6]+tmp[5086]*kernel[7]+tmp[5087]*kernel[8];
				ans[4987]<=tmp[4886]*kernel[0]+tmp[4887]*kernel[1]+tmp[4888]*kernel[2]+tmp[4986]*kernel[3]+tmp[4987]*kernel[4]+tmp[4988]*kernel[5]+tmp[5086]*kernel[6]+tmp[5087]*kernel[7]+tmp[5088]*kernel[8];
				ans[4988]<=tmp[4887]*kernel[0]+tmp[4888]*kernel[1]+tmp[4889]*kernel[2]+tmp[4987]*kernel[3]+tmp[4988]*kernel[4]+tmp[4989]*kernel[5]+tmp[5087]*kernel[6]+tmp[5088]*kernel[7]+tmp[5089]*kernel[8];
				ans[4989]<=tmp[4888]*kernel[0]+tmp[4889]*kernel[1]+tmp[4890]*kernel[2]+tmp[4988]*kernel[3]+tmp[4989]*kernel[4]+tmp[4990]*kernel[5]+tmp[5088]*kernel[6]+tmp[5089]*kernel[7]+tmp[5090]*kernel[8];
				ans[4990]<=tmp[4889]*kernel[0]+tmp[4890]*kernel[1]+tmp[4891]*kernel[2]+tmp[4989]*kernel[3]+tmp[4990]*kernel[4]+tmp[4991]*kernel[5]+tmp[5089]*kernel[6]+tmp[5090]*kernel[7]+tmp[5091]*kernel[8];
				ans[4991]<=tmp[4890]*kernel[0]+tmp[4891]*kernel[1]+tmp[4892]*kernel[2]+tmp[4990]*kernel[3]+tmp[4991]*kernel[4]+tmp[4992]*kernel[5]+tmp[5090]*kernel[6]+tmp[5091]*kernel[7]+tmp[5092]*kernel[8];
				ans[4992]<=tmp[4891]*kernel[0]+tmp[4892]*kernel[1]+tmp[4893]*kernel[2]+tmp[4991]*kernel[3]+tmp[4992]*kernel[4]+tmp[4993]*kernel[5]+tmp[5091]*kernel[6]+tmp[5092]*kernel[7]+tmp[5093]*kernel[8];
				ans[4993]<=tmp[4892]*kernel[0]+tmp[4893]*kernel[1]+tmp[4894]*kernel[2]+tmp[4992]*kernel[3]+tmp[4993]*kernel[4]+tmp[4994]*kernel[5]+tmp[5092]*kernel[6]+tmp[5093]*kernel[7]+tmp[5094]*kernel[8];
				ans[4994]<=tmp[4893]*kernel[0]+tmp[4894]*kernel[1]+tmp[4895]*kernel[2]+tmp[4993]*kernel[3]+tmp[4994]*kernel[4]+tmp[4995]*kernel[5]+tmp[5093]*kernel[6]+tmp[5094]*kernel[7]+tmp[5095]*kernel[8];
				ans[4995]<=tmp[4894]*kernel[0]+tmp[4895]*kernel[1]+tmp[4896]*kernel[2]+tmp[4994]*kernel[3]+tmp[4995]*kernel[4]+tmp[4996]*kernel[5]+tmp[5094]*kernel[6]+tmp[5095]*kernel[7]+tmp[5096]*kernel[8];
				ans[4996]<=tmp[4895]*kernel[0]+tmp[4896]*kernel[1]+tmp[4897]*kernel[2]+tmp[4995]*kernel[3]+tmp[4996]*kernel[4]+tmp[4997]*kernel[5]+tmp[5095]*kernel[6]+tmp[5096]*kernel[7]+tmp[5097]*kernel[8];
				ans[4997]<=tmp[4896]*kernel[0]+tmp[4897]*kernel[1]+tmp[4898]*kernel[2]+tmp[4996]*kernel[3]+tmp[4997]*kernel[4]+tmp[4998]*kernel[5]+tmp[5096]*kernel[6]+tmp[5097]*kernel[7]+tmp[5098]*kernel[8];
				ans[4998]<=tmp[4897]*kernel[0]+tmp[4898]*kernel[1]+tmp[4899]*kernel[2]+tmp[4997]*kernel[3]+tmp[4998]*kernel[4]+tmp[4999]*kernel[5]+tmp[5097]*kernel[6]+tmp[5098]*kernel[7]+tmp[5099]*kernel[8];
				ans[4999]<=tmp[4898]*kernel[0]+tmp[4899]*kernel[1]+tmp[4998]*kernel[3]+tmp[4999]*kernel[4]+tmp[5098]*kernel[6]+tmp[5099]*kernel[7];
				ans[5000]<=tmp[4900]*kernel[1]+tmp[4901]*kernel[2]+tmp[5000]*kernel[4]+tmp[5001]*kernel[5]+tmp[5100]*kernel[7]+tmp[5101]*kernel[8];
				ans[5001]<=tmp[4900]*kernel[0]+tmp[4901]*kernel[1]+tmp[4902]*kernel[2]+tmp[5000]*kernel[3]+tmp[5001]*kernel[4]+tmp[5002]*kernel[5]+tmp[5100]*kernel[6]+tmp[5101]*kernel[7]+tmp[5102]*kernel[8];
				ans[5002]<=tmp[4901]*kernel[0]+tmp[4902]*kernel[1]+tmp[4903]*kernel[2]+tmp[5001]*kernel[3]+tmp[5002]*kernel[4]+tmp[5003]*kernel[5]+tmp[5101]*kernel[6]+tmp[5102]*kernel[7]+tmp[5103]*kernel[8];
				ans[5003]<=tmp[4902]*kernel[0]+tmp[4903]*kernel[1]+tmp[4904]*kernel[2]+tmp[5002]*kernel[3]+tmp[5003]*kernel[4]+tmp[5004]*kernel[5]+tmp[5102]*kernel[6]+tmp[5103]*kernel[7]+tmp[5104]*kernel[8];
				ans[5004]<=tmp[4903]*kernel[0]+tmp[4904]*kernel[1]+tmp[4905]*kernel[2]+tmp[5003]*kernel[3]+tmp[5004]*kernel[4]+tmp[5005]*kernel[5]+tmp[5103]*kernel[6]+tmp[5104]*kernel[7]+tmp[5105]*kernel[8];
				ans[5005]<=tmp[4904]*kernel[0]+tmp[4905]*kernel[1]+tmp[4906]*kernel[2]+tmp[5004]*kernel[3]+tmp[5005]*kernel[4]+tmp[5006]*kernel[5]+tmp[5104]*kernel[6]+tmp[5105]*kernel[7]+tmp[5106]*kernel[8];
				ans[5006]<=tmp[4905]*kernel[0]+tmp[4906]*kernel[1]+tmp[4907]*kernel[2]+tmp[5005]*kernel[3]+tmp[5006]*kernel[4]+tmp[5007]*kernel[5]+tmp[5105]*kernel[6]+tmp[5106]*kernel[7]+tmp[5107]*kernel[8];
				ans[5007]<=tmp[4906]*kernel[0]+tmp[4907]*kernel[1]+tmp[4908]*kernel[2]+tmp[5006]*kernel[3]+tmp[5007]*kernel[4]+tmp[5008]*kernel[5]+tmp[5106]*kernel[6]+tmp[5107]*kernel[7]+tmp[5108]*kernel[8];
				ans[5008]<=tmp[4907]*kernel[0]+tmp[4908]*kernel[1]+tmp[4909]*kernel[2]+tmp[5007]*kernel[3]+tmp[5008]*kernel[4]+tmp[5009]*kernel[5]+tmp[5107]*kernel[6]+tmp[5108]*kernel[7]+tmp[5109]*kernel[8];
				ans[5009]<=tmp[4908]*kernel[0]+tmp[4909]*kernel[1]+tmp[4910]*kernel[2]+tmp[5008]*kernel[3]+tmp[5009]*kernel[4]+tmp[5010]*kernel[5]+tmp[5108]*kernel[6]+tmp[5109]*kernel[7]+tmp[5110]*kernel[8];
				ans[5010]<=tmp[4909]*kernel[0]+tmp[4910]*kernel[1]+tmp[4911]*kernel[2]+tmp[5009]*kernel[3]+tmp[5010]*kernel[4]+tmp[5011]*kernel[5]+tmp[5109]*kernel[6]+tmp[5110]*kernel[7]+tmp[5111]*kernel[8];
				ans[5011]<=tmp[4910]*kernel[0]+tmp[4911]*kernel[1]+tmp[4912]*kernel[2]+tmp[5010]*kernel[3]+tmp[5011]*kernel[4]+tmp[5012]*kernel[5]+tmp[5110]*kernel[6]+tmp[5111]*kernel[7]+tmp[5112]*kernel[8];
				ans[5012]<=tmp[4911]*kernel[0]+tmp[4912]*kernel[1]+tmp[4913]*kernel[2]+tmp[5011]*kernel[3]+tmp[5012]*kernel[4]+tmp[5013]*kernel[5]+tmp[5111]*kernel[6]+tmp[5112]*kernel[7]+tmp[5113]*kernel[8];
				ans[5013]<=tmp[4912]*kernel[0]+tmp[4913]*kernel[1]+tmp[4914]*kernel[2]+tmp[5012]*kernel[3]+tmp[5013]*kernel[4]+tmp[5014]*kernel[5]+tmp[5112]*kernel[6]+tmp[5113]*kernel[7]+tmp[5114]*kernel[8];
				ans[5014]<=tmp[4913]*kernel[0]+tmp[4914]*kernel[1]+tmp[4915]*kernel[2]+tmp[5013]*kernel[3]+tmp[5014]*kernel[4]+tmp[5015]*kernel[5]+tmp[5113]*kernel[6]+tmp[5114]*kernel[7]+tmp[5115]*kernel[8];
				ans[5015]<=tmp[4914]*kernel[0]+tmp[4915]*kernel[1]+tmp[4916]*kernel[2]+tmp[5014]*kernel[3]+tmp[5015]*kernel[4]+tmp[5016]*kernel[5]+tmp[5114]*kernel[6]+tmp[5115]*kernel[7]+tmp[5116]*kernel[8];
				ans[5016]<=tmp[4915]*kernel[0]+tmp[4916]*kernel[1]+tmp[4917]*kernel[2]+tmp[5015]*kernel[3]+tmp[5016]*kernel[4]+tmp[5017]*kernel[5]+tmp[5115]*kernel[6]+tmp[5116]*kernel[7]+tmp[5117]*kernel[8];
				ans[5017]<=tmp[4916]*kernel[0]+tmp[4917]*kernel[1]+tmp[4918]*kernel[2]+tmp[5016]*kernel[3]+tmp[5017]*kernel[4]+tmp[5018]*kernel[5]+tmp[5116]*kernel[6]+tmp[5117]*kernel[7]+tmp[5118]*kernel[8];
				ans[5018]<=tmp[4917]*kernel[0]+tmp[4918]*kernel[1]+tmp[4919]*kernel[2]+tmp[5017]*kernel[3]+tmp[5018]*kernel[4]+tmp[5019]*kernel[5]+tmp[5117]*kernel[6]+tmp[5118]*kernel[7]+tmp[5119]*kernel[8];
				ans[5019]<=tmp[4918]*kernel[0]+tmp[4919]*kernel[1]+tmp[4920]*kernel[2]+tmp[5018]*kernel[3]+tmp[5019]*kernel[4]+tmp[5020]*kernel[5]+tmp[5118]*kernel[6]+tmp[5119]*kernel[7]+tmp[5120]*kernel[8];
				ans[5020]<=tmp[4919]*kernel[0]+tmp[4920]*kernel[1]+tmp[4921]*kernel[2]+tmp[5019]*kernel[3]+tmp[5020]*kernel[4]+tmp[5021]*kernel[5]+tmp[5119]*kernel[6]+tmp[5120]*kernel[7]+tmp[5121]*kernel[8];
				ans[5021]<=tmp[4920]*kernel[0]+tmp[4921]*kernel[1]+tmp[4922]*kernel[2]+tmp[5020]*kernel[3]+tmp[5021]*kernel[4]+tmp[5022]*kernel[5]+tmp[5120]*kernel[6]+tmp[5121]*kernel[7]+tmp[5122]*kernel[8];
				ans[5022]<=tmp[4921]*kernel[0]+tmp[4922]*kernel[1]+tmp[4923]*kernel[2]+tmp[5021]*kernel[3]+tmp[5022]*kernel[4]+tmp[5023]*kernel[5]+tmp[5121]*kernel[6]+tmp[5122]*kernel[7]+tmp[5123]*kernel[8];
				ans[5023]<=tmp[4922]*kernel[0]+tmp[4923]*kernel[1]+tmp[4924]*kernel[2]+tmp[5022]*kernel[3]+tmp[5023]*kernel[4]+tmp[5024]*kernel[5]+tmp[5122]*kernel[6]+tmp[5123]*kernel[7]+tmp[5124]*kernel[8];
				ans[5024]<=tmp[4923]*kernel[0]+tmp[4924]*kernel[1]+tmp[4925]*kernel[2]+tmp[5023]*kernel[3]+tmp[5024]*kernel[4]+tmp[5025]*kernel[5]+tmp[5123]*kernel[6]+tmp[5124]*kernel[7]+tmp[5125]*kernel[8];
				ans[5025]<=tmp[4924]*kernel[0]+tmp[4925]*kernel[1]+tmp[4926]*kernel[2]+tmp[5024]*kernel[3]+tmp[5025]*kernel[4]+tmp[5026]*kernel[5]+tmp[5124]*kernel[6]+tmp[5125]*kernel[7]+tmp[5126]*kernel[8];
				ans[5026]<=tmp[4925]*kernel[0]+tmp[4926]*kernel[1]+tmp[4927]*kernel[2]+tmp[5025]*kernel[3]+tmp[5026]*kernel[4]+tmp[5027]*kernel[5]+tmp[5125]*kernel[6]+tmp[5126]*kernel[7]+tmp[5127]*kernel[8];
				ans[5027]<=tmp[4926]*kernel[0]+tmp[4927]*kernel[1]+tmp[4928]*kernel[2]+tmp[5026]*kernel[3]+tmp[5027]*kernel[4]+tmp[5028]*kernel[5]+tmp[5126]*kernel[6]+tmp[5127]*kernel[7]+tmp[5128]*kernel[8];
				ans[5028]<=tmp[4927]*kernel[0]+tmp[4928]*kernel[1]+tmp[4929]*kernel[2]+tmp[5027]*kernel[3]+tmp[5028]*kernel[4]+tmp[5029]*kernel[5]+tmp[5127]*kernel[6]+tmp[5128]*kernel[7]+tmp[5129]*kernel[8];
				ans[5029]<=tmp[4928]*kernel[0]+tmp[4929]*kernel[1]+tmp[4930]*kernel[2]+tmp[5028]*kernel[3]+tmp[5029]*kernel[4]+tmp[5030]*kernel[5]+tmp[5128]*kernel[6]+tmp[5129]*kernel[7]+tmp[5130]*kernel[8];
				ans[5030]<=tmp[4929]*kernel[0]+tmp[4930]*kernel[1]+tmp[4931]*kernel[2]+tmp[5029]*kernel[3]+tmp[5030]*kernel[4]+tmp[5031]*kernel[5]+tmp[5129]*kernel[6]+tmp[5130]*kernel[7]+tmp[5131]*kernel[8];
				ans[5031]<=tmp[4930]*kernel[0]+tmp[4931]*kernel[1]+tmp[4932]*kernel[2]+tmp[5030]*kernel[3]+tmp[5031]*kernel[4]+tmp[5032]*kernel[5]+tmp[5130]*kernel[6]+tmp[5131]*kernel[7]+tmp[5132]*kernel[8];
				ans[5032]<=tmp[4931]*kernel[0]+tmp[4932]*kernel[1]+tmp[4933]*kernel[2]+tmp[5031]*kernel[3]+tmp[5032]*kernel[4]+tmp[5033]*kernel[5]+tmp[5131]*kernel[6]+tmp[5132]*kernel[7]+tmp[5133]*kernel[8];
				ans[5033]<=tmp[4932]*kernel[0]+tmp[4933]*kernel[1]+tmp[4934]*kernel[2]+tmp[5032]*kernel[3]+tmp[5033]*kernel[4]+tmp[5034]*kernel[5]+tmp[5132]*kernel[6]+tmp[5133]*kernel[7]+tmp[5134]*kernel[8];
				ans[5034]<=tmp[4933]*kernel[0]+tmp[4934]*kernel[1]+tmp[4935]*kernel[2]+tmp[5033]*kernel[3]+tmp[5034]*kernel[4]+tmp[5035]*kernel[5]+tmp[5133]*kernel[6]+tmp[5134]*kernel[7]+tmp[5135]*kernel[8];
				ans[5035]<=tmp[4934]*kernel[0]+tmp[4935]*kernel[1]+tmp[4936]*kernel[2]+tmp[5034]*kernel[3]+tmp[5035]*kernel[4]+tmp[5036]*kernel[5]+tmp[5134]*kernel[6]+tmp[5135]*kernel[7]+tmp[5136]*kernel[8];
				ans[5036]<=tmp[4935]*kernel[0]+tmp[4936]*kernel[1]+tmp[4937]*kernel[2]+tmp[5035]*kernel[3]+tmp[5036]*kernel[4]+tmp[5037]*kernel[5]+tmp[5135]*kernel[6]+tmp[5136]*kernel[7]+tmp[5137]*kernel[8];
				ans[5037]<=tmp[4936]*kernel[0]+tmp[4937]*kernel[1]+tmp[4938]*kernel[2]+tmp[5036]*kernel[3]+tmp[5037]*kernel[4]+tmp[5038]*kernel[5]+tmp[5136]*kernel[6]+tmp[5137]*kernel[7]+tmp[5138]*kernel[8];
				ans[5038]<=tmp[4937]*kernel[0]+tmp[4938]*kernel[1]+tmp[4939]*kernel[2]+tmp[5037]*kernel[3]+tmp[5038]*kernel[4]+tmp[5039]*kernel[5]+tmp[5137]*kernel[6]+tmp[5138]*kernel[7]+tmp[5139]*kernel[8];
				ans[5039]<=tmp[4938]*kernel[0]+tmp[4939]*kernel[1]+tmp[4940]*kernel[2]+tmp[5038]*kernel[3]+tmp[5039]*kernel[4]+tmp[5040]*kernel[5]+tmp[5138]*kernel[6]+tmp[5139]*kernel[7]+tmp[5140]*kernel[8];
				ans[5040]<=tmp[4939]*kernel[0]+tmp[4940]*kernel[1]+tmp[4941]*kernel[2]+tmp[5039]*kernel[3]+tmp[5040]*kernel[4]+tmp[5041]*kernel[5]+tmp[5139]*kernel[6]+tmp[5140]*kernel[7]+tmp[5141]*kernel[8];
				ans[5041]<=tmp[4940]*kernel[0]+tmp[4941]*kernel[1]+tmp[4942]*kernel[2]+tmp[5040]*kernel[3]+tmp[5041]*kernel[4]+tmp[5042]*kernel[5]+tmp[5140]*kernel[6]+tmp[5141]*kernel[7]+tmp[5142]*kernel[8];
				ans[5042]<=tmp[4941]*kernel[0]+tmp[4942]*kernel[1]+tmp[4943]*kernel[2]+tmp[5041]*kernel[3]+tmp[5042]*kernel[4]+tmp[5043]*kernel[5]+tmp[5141]*kernel[6]+tmp[5142]*kernel[7]+tmp[5143]*kernel[8];
				ans[5043]<=tmp[4942]*kernel[0]+tmp[4943]*kernel[1]+tmp[4944]*kernel[2]+tmp[5042]*kernel[3]+tmp[5043]*kernel[4]+tmp[5044]*kernel[5]+tmp[5142]*kernel[6]+tmp[5143]*kernel[7]+tmp[5144]*kernel[8];
				ans[5044]<=tmp[4943]*kernel[0]+tmp[4944]*kernel[1]+tmp[4945]*kernel[2]+tmp[5043]*kernel[3]+tmp[5044]*kernel[4]+tmp[5045]*kernel[5]+tmp[5143]*kernel[6]+tmp[5144]*kernel[7]+tmp[5145]*kernel[8];
				ans[5045]<=tmp[4944]*kernel[0]+tmp[4945]*kernel[1]+tmp[4946]*kernel[2]+tmp[5044]*kernel[3]+tmp[5045]*kernel[4]+tmp[5046]*kernel[5]+tmp[5144]*kernel[6]+tmp[5145]*kernel[7]+tmp[5146]*kernel[8];
				ans[5046]<=tmp[4945]*kernel[0]+tmp[4946]*kernel[1]+tmp[4947]*kernel[2]+tmp[5045]*kernel[3]+tmp[5046]*kernel[4]+tmp[5047]*kernel[5]+tmp[5145]*kernel[6]+tmp[5146]*kernel[7]+tmp[5147]*kernel[8];
				ans[5047]<=tmp[4946]*kernel[0]+tmp[4947]*kernel[1]+tmp[4948]*kernel[2]+tmp[5046]*kernel[3]+tmp[5047]*kernel[4]+tmp[5048]*kernel[5]+tmp[5146]*kernel[6]+tmp[5147]*kernel[7]+tmp[5148]*kernel[8];
				ans[5048]<=tmp[4947]*kernel[0]+tmp[4948]*kernel[1]+tmp[4949]*kernel[2]+tmp[5047]*kernel[3]+tmp[5048]*kernel[4]+tmp[5049]*kernel[5]+tmp[5147]*kernel[6]+tmp[5148]*kernel[7]+tmp[5149]*kernel[8];
				ans[5049]<=tmp[4948]*kernel[0]+tmp[4949]*kernel[1]+tmp[4950]*kernel[2]+tmp[5048]*kernel[3]+tmp[5049]*kernel[4]+tmp[5050]*kernel[5]+tmp[5148]*kernel[6]+tmp[5149]*kernel[7]+tmp[5150]*kernel[8];
				ans[5050]<=tmp[4949]*kernel[0]+tmp[4950]*kernel[1]+tmp[4951]*kernel[2]+tmp[5049]*kernel[3]+tmp[5050]*kernel[4]+tmp[5051]*kernel[5]+tmp[5149]*kernel[6]+tmp[5150]*kernel[7]+tmp[5151]*kernel[8];
				ans[5051]<=tmp[4950]*kernel[0]+tmp[4951]*kernel[1]+tmp[4952]*kernel[2]+tmp[5050]*kernel[3]+tmp[5051]*kernel[4]+tmp[5052]*kernel[5]+tmp[5150]*kernel[6]+tmp[5151]*kernel[7]+tmp[5152]*kernel[8];
				ans[5052]<=tmp[4951]*kernel[0]+tmp[4952]*kernel[1]+tmp[4953]*kernel[2]+tmp[5051]*kernel[3]+tmp[5052]*kernel[4]+tmp[5053]*kernel[5]+tmp[5151]*kernel[6]+tmp[5152]*kernel[7]+tmp[5153]*kernel[8];
				ans[5053]<=tmp[4952]*kernel[0]+tmp[4953]*kernel[1]+tmp[4954]*kernel[2]+tmp[5052]*kernel[3]+tmp[5053]*kernel[4]+tmp[5054]*kernel[5]+tmp[5152]*kernel[6]+tmp[5153]*kernel[7]+tmp[5154]*kernel[8];
				ans[5054]<=tmp[4953]*kernel[0]+tmp[4954]*kernel[1]+tmp[4955]*kernel[2]+tmp[5053]*kernel[3]+tmp[5054]*kernel[4]+tmp[5055]*kernel[5]+tmp[5153]*kernel[6]+tmp[5154]*kernel[7]+tmp[5155]*kernel[8];
				ans[5055]<=tmp[4954]*kernel[0]+tmp[4955]*kernel[1]+tmp[4956]*kernel[2]+tmp[5054]*kernel[3]+tmp[5055]*kernel[4]+tmp[5056]*kernel[5]+tmp[5154]*kernel[6]+tmp[5155]*kernel[7]+tmp[5156]*kernel[8];
				ans[5056]<=tmp[4955]*kernel[0]+tmp[4956]*kernel[1]+tmp[4957]*kernel[2]+tmp[5055]*kernel[3]+tmp[5056]*kernel[4]+tmp[5057]*kernel[5]+tmp[5155]*kernel[6]+tmp[5156]*kernel[7]+tmp[5157]*kernel[8];
				ans[5057]<=tmp[4956]*kernel[0]+tmp[4957]*kernel[1]+tmp[4958]*kernel[2]+tmp[5056]*kernel[3]+tmp[5057]*kernel[4]+tmp[5058]*kernel[5]+tmp[5156]*kernel[6]+tmp[5157]*kernel[7]+tmp[5158]*kernel[8];
				ans[5058]<=tmp[4957]*kernel[0]+tmp[4958]*kernel[1]+tmp[4959]*kernel[2]+tmp[5057]*kernel[3]+tmp[5058]*kernel[4]+tmp[5059]*kernel[5]+tmp[5157]*kernel[6]+tmp[5158]*kernel[7]+tmp[5159]*kernel[8];
				ans[5059]<=tmp[4958]*kernel[0]+tmp[4959]*kernel[1]+tmp[4960]*kernel[2]+tmp[5058]*kernel[3]+tmp[5059]*kernel[4]+tmp[5060]*kernel[5]+tmp[5158]*kernel[6]+tmp[5159]*kernel[7]+tmp[5160]*kernel[8];
				ans[5060]<=tmp[4959]*kernel[0]+tmp[4960]*kernel[1]+tmp[4961]*kernel[2]+tmp[5059]*kernel[3]+tmp[5060]*kernel[4]+tmp[5061]*kernel[5]+tmp[5159]*kernel[6]+tmp[5160]*kernel[7]+tmp[5161]*kernel[8];
				ans[5061]<=tmp[4960]*kernel[0]+tmp[4961]*kernel[1]+tmp[4962]*kernel[2]+tmp[5060]*kernel[3]+tmp[5061]*kernel[4]+tmp[5062]*kernel[5]+tmp[5160]*kernel[6]+tmp[5161]*kernel[7]+tmp[5162]*kernel[8];
				ans[5062]<=tmp[4961]*kernel[0]+tmp[4962]*kernel[1]+tmp[4963]*kernel[2]+tmp[5061]*kernel[3]+tmp[5062]*kernel[4]+tmp[5063]*kernel[5]+tmp[5161]*kernel[6]+tmp[5162]*kernel[7]+tmp[5163]*kernel[8];
				ans[5063]<=tmp[4962]*kernel[0]+tmp[4963]*kernel[1]+tmp[4964]*kernel[2]+tmp[5062]*kernel[3]+tmp[5063]*kernel[4]+tmp[5064]*kernel[5]+tmp[5162]*kernel[6]+tmp[5163]*kernel[7]+tmp[5164]*kernel[8];
				ans[5064]<=tmp[4963]*kernel[0]+tmp[4964]*kernel[1]+tmp[4965]*kernel[2]+tmp[5063]*kernel[3]+tmp[5064]*kernel[4]+tmp[5065]*kernel[5]+tmp[5163]*kernel[6]+tmp[5164]*kernel[7]+tmp[5165]*kernel[8];
				ans[5065]<=tmp[4964]*kernel[0]+tmp[4965]*kernel[1]+tmp[4966]*kernel[2]+tmp[5064]*kernel[3]+tmp[5065]*kernel[4]+tmp[5066]*kernel[5]+tmp[5164]*kernel[6]+tmp[5165]*kernel[7]+tmp[5166]*kernel[8];
				ans[5066]<=tmp[4965]*kernel[0]+tmp[4966]*kernel[1]+tmp[4967]*kernel[2]+tmp[5065]*kernel[3]+tmp[5066]*kernel[4]+tmp[5067]*kernel[5]+tmp[5165]*kernel[6]+tmp[5166]*kernel[7]+tmp[5167]*kernel[8];
				ans[5067]<=tmp[4966]*kernel[0]+tmp[4967]*kernel[1]+tmp[4968]*kernel[2]+tmp[5066]*kernel[3]+tmp[5067]*kernel[4]+tmp[5068]*kernel[5]+tmp[5166]*kernel[6]+tmp[5167]*kernel[7]+tmp[5168]*kernel[8];
				ans[5068]<=tmp[4967]*kernel[0]+tmp[4968]*kernel[1]+tmp[4969]*kernel[2]+tmp[5067]*kernel[3]+tmp[5068]*kernel[4]+tmp[5069]*kernel[5]+tmp[5167]*kernel[6]+tmp[5168]*kernel[7]+tmp[5169]*kernel[8];
				ans[5069]<=tmp[4968]*kernel[0]+tmp[4969]*kernel[1]+tmp[4970]*kernel[2]+tmp[5068]*kernel[3]+tmp[5069]*kernel[4]+tmp[5070]*kernel[5]+tmp[5168]*kernel[6]+tmp[5169]*kernel[7]+tmp[5170]*kernel[8];
				ans[5070]<=tmp[4969]*kernel[0]+tmp[4970]*kernel[1]+tmp[4971]*kernel[2]+tmp[5069]*kernel[3]+tmp[5070]*kernel[4]+tmp[5071]*kernel[5]+tmp[5169]*kernel[6]+tmp[5170]*kernel[7]+tmp[5171]*kernel[8];
				ans[5071]<=tmp[4970]*kernel[0]+tmp[4971]*kernel[1]+tmp[4972]*kernel[2]+tmp[5070]*kernel[3]+tmp[5071]*kernel[4]+tmp[5072]*kernel[5]+tmp[5170]*kernel[6]+tmp[5171]*kernel[7]+tmp[5172]*kernel[8];
				ans[5072]<=tmp[4971]*kernel[0]+tmp[4972]*kernel[1]+tmp[4973]*kernel[2]+tmp[5071]*kernel[3]+tmp[5072]*kernel[4]+tmp[5073]*kernel[5]+tmp[5171]*kernel[6]+tmp[5172]*kernel[7]+tmp[5173]*kernel[8];
				ans[5073]<=tmp[4972]*kernel[0]+tmp[4973]*kernel[1]+tmp[4974]*kernel[2]+tmp[5072]*kernel[3]+tmp[5073]*kernel[4]+tmp[5074]*kernel[5]+tmp[5172]*kernel[6]+tmp[5173]*kernel[7]+tmp[5174]*kernel[8];
				ans[5074]<=tmp[4973]*kernel[0]+tmp[4974]*kernel[1]+tmp[4975]*kernel[2]+tmp[5073]*kernel[3]+tmp[5074]*kernel[4]+tmp[5075]*kernel[5]+tmp[5173]*kernel[6]+tmp[5174]*kernel[7]+tmp[5175]*kernel[8];
				ans[5075]<=tmp[4974]*kernel[0]+tmp[4975]*kernel[1]+tmp[4976]*kernel[2]+tmp[5074]*kernel[3]+tmp[5075]*kernel[4]+tmp[5076]*kernel[5]+tmp[5174]*kernel[6]+tmp[5175]*kernel[7]+tmp[5176]*kernel[8];
				ans[5076]<=tmp[4975]*kernel[0]+tmp[4976]*kernel[1]+tmp[4977]*kernel[2]+tmp[5075]*kernel[3]+tmp[5076]*kernel[4]+tmp[5077]*kernel[5]+tmp[5175]*kernel[6]+tmp[5176]*kernel[7]+tmp[5177]*kernel[8];
				ans[5077]<=tmp[4976]*kernel[0]+tmp[4977]*kernel[1]+tmp[4978]*kernel[2]+tmp[5076]*kernel[3]+tmp[5077]*kernel[4]+tmp[5078]*kernel[5]+tmp[5176]*kernel[6]+tmp[5177]*kernel[7]+tmp[5178]*kernel[8];
				ans[5078]<=tmp[4977]*kernel[0]+tmp[4978]*kernel[1]+tmp[4979]*kernel[2]+tmp[5077]*kernel[3]+tmp[5078]*kernel[4]+tmp[5079]*kernel[5]+tmp[5177]*kernel[6]+tmp[5178]*kernel[7]+tmp[5179]*kernel[8];
				ans[5079]<=tmp[4978]*kernel[0]+tmp[4979]*kernel[1]+tmp[4980]*kernel[2]+tmp[5078]*kernel[3]+tmp[5079]*kernel[4]+tmp[5080]*kernel[5]+tmp[5178]*kernel[6]+tmp[5179]*kernel[7]+tmp[5180]*kernel[8];
				ans[5080]<=tmp[4979]*kernel[0]+tmp[4980]*kernel[1]+tmp[4981]*kernel[2]+tmp[5079]*kernel[3]+tmp[5080]*kernel[4]+tmp[5081]*kernel[5]+tmp[5179]*kernel[6]+tmp[5180]*kernel[7]+tmp[5181]*kernel[8];
				ans[5081]<=tmp[4980]*kernel[0]+tmp[4981]*kernel[1]+tmp[4982]*kernel[2]+tmp[5080]*kernel[3]+tmp[5081]*kernel[4]+tmp[5082]*kernel[5]+tmp[5180]*kernel[6]+tmp[5181]*kernel[7]+tmp[5182]*kernel[8];
				ans[5082]<=tmp[4981]*kernel[0]+tmp[4982]*kernel[1]+tmp[4983]*kernel[2]+tmp[5081]*kernel[3]+tmp[5082]*kernel[4]+tmp[5083]*kernel[5]+tmp[5181]*kernel[6]+tmp[5182]*kernel[7]+tmp[5183]*kernel[8];
				ans[5083]<=tmp[4982]*kernel[0]+tmp[4983]*kernel[1]+tmp[4984]*kernel[2]+tmp[5082]*kernel[3]+tmp[5083]*kernel[4]+tmp[5084]*kernel[5]+tmp[5182]*kernel[6]+tmp[5183]*kernel[7]+tmp[5184]*kernel[8];
				ans[5084]<=tmp[4983]*kernel[0]+tmp[4984]*kernel[1]+tmp[4985]*kernel[2]+tmp[5083]*kernel[3]+tmp[5084]*kernel[4]+tmp[5085]*kernel[5]+tmp[5183]*kernel[6]+tmp[5184]*kernel[7]+tmp[5185]*kernel[8];
				ans[5085]<=tmp[4984]*kernel[0]+tmp[4985]*kernel[1]+tmp[4986]*kernel[2]+tmp[5084]*kernel[3]+tmp[5085]*kernel[4]+tmp[5086]*kernel[5]+tmp[5184]*kernel[6]+tmp[5185]*kernel[7]+tmp[5186]*kernel[8];
				ans[5086]<=tmp[4985]*kernel[0]+tmp[4986]*kernel[1]+tmp[4987]*kernel[2]+tmp[5085]*kernel[3]+tmp[5086]*kernel[4]+tmp[5087]*kernel[5]+tmp[5185]*kernel[6]+tmp[5186]*kernel[7]+tmp[5187]*kernel[8];
				ans[5087]<=tmp[4986]*kernel[0]+tmp[4987]*kernel[1]+tmp[4988]*kernel[2]+tmp[5086]*kernel[3]+tmp[5087]*kernel[4]+tmp[5088]*kernel[5]+tmp[5186]*kernel[6]+tmp[5187]*kernel[7]+tmp[5188]*kernel[8];
				ans[5088]<=tmp[4987]*kernel[0]+tmp[4988]*kernel[1]+tmp[4989]*kernel[2]+tmp[5087]*kernel[3]+tmp[5088]*kernel[4]+tmp[5089]*kernel[5]+tmp[5187]*kernel[6]+tmp[5188]*kernel[7]+tmp[5189]*kernel[8];
				ans[5089]<=tmp[4988]*kernel[0]+tmp[4989]*kernel[1]+tmp[4990]*kernel[2]+tmp[5088]*kernel[3]+tmp[5089]*kernel[4]+tmp[5090]*kernel[5]+tmp[5188]*kernel[6]+tmp[5189]*kernel[7]+tmp[5190]*kernel[8];
				ans[5090]<=tmp[4989]*kernel[0]+tmp[4990]*kernel[1]+tmp[4991]*kernel[2]+tmp[5089]*kernel[3]+tmp[5090]*kernel[4]+tmp[5091]*kernel[5]+tmp[5189]*kernel[6]+tmp[5190]*kernel[7]+tmp[5191]*kernel[8];
				ans[5091]<=tmp[4990]*kernel[0]+tmp[4991]*kernel[1]+tmp[4992]*kernel[2]+tmp[5090]*kernel[3]+tmp[5091]*kernel[4]+tmp[5092]*kernel[5]+tmp[5190]*kernel[6]+tmp[5191]*kernel[7]+tmp[5192]*kernel[8];
				ans[5092]<=tmp[4991]*kernel[0]+tmp[4992]*kernel[1]+tmp[4993]*kernel[2]+tmp[5091]*kernel[3]+tmp[5092]*kernel[4]+tmp[5093]*kernel[5]+tmp[5191]*kernel[6]+tmp[5192]*kernel[7]+tmp[5193]*kernel[8];
				ans[5093]<=tmp[4992]*kernel[0]+tmp[4993]*kernel[1]+tmp[4994]*kernel[2]+tmp[5092]*kernel[3]+tmp[5093]*kernel[4]+tmp[5094]*kernel[5]+tmp[5192]*kernel[6]+tmp[5193]*kernel[7]+tmp[5194]*kernel[8];
				ans[5094]<=tmp[4993]*kernel[0]+tmp[4994]*kernel[1]+tmp[4995]*kernel[2]+tmp[5093]*kernel[3]+tmp[5094]*kernel[4]+tmp[5095]*kernel[5]+tmp[5193]*kernel[6]+tmp[5194]*kernel[7]+tmp[5195]*kernel[8];
				ans[5095]<=tmp[4994]*kernel[0]+tmp[4995]*kernel[1]+tmp[4996]*kernel[2]+tmp[5094]*kernel[3]+tmp[5095]*kernel[4]+tmp[5096]*kernel[5]+tmp[5194]*kernel[6]+tmp[5195]*kernel[7]+tmp[5196]*kernel[8];
				ans[5096]<=tmp[4995]*kernel[0]+tmp[4996]*kernel[1]+tmp[4997]*kernel[2]+tmp[5095]*kernel[3]+tmp[5096]*kernel[4]+tmp[5097]*kernel[5]+tmp[5195]*kernel[6]+tmp[5196]*kernel[7]+tmp[5197]*kernel[8];
				ans[5097]<=tmp[4996]*kernel[0]+tmp[4997]*kernel[1]+tmp[4998]*kernel[2]+tmp[5096]*kernel[3]+tmp[5097]*kernel[4]+tmp[5098]*kernel[5]+tmp[5196]*kernel[6]+tmp[5197]*kernel[7]+tmp[5198]*kernel[8];
				ans[5098]<=tmp[4997]*kernel[0]+tmp[4998]*kernel[1]+tmp[4999]*kernel[2]+tmp[5097]*kernel[3]+tmp[5098]*kernel[4]+tmp[5099]*kernel[5]+tmp[5197]*kernel[6]+tmp[5198]*kernel[7]+tmp[5199]*kernel[8];
				ans[5099]<=tmp[4998]*kernel[0]+tmp[4999]*kernel[1]+tmp[5098]*kernel[3]+tmp[5099]*kernel[4]+tmp[5198]*kernel[6]+tmp[5199]*kernel[7];
				ans[5100]<=tmp[5000]*kernel[1]+tmp[5001]*kernel[2]+tmp[5100]*kernel[4]+tmp[5101]*kernel[5]+tmp[5200]*kernel[7]+tmp[5201]*kernel[8];
				ans[5101]<=tmp[5000]*kernel[0]+tmp[5001]*kernel[1]+tmp[5002]*kernel[2]+tmp[5100]*kernel[3]+tmp[5101]*kernel[4]+tmp[5102]*kernel[5]+tmp[5200]*kernel[6]+tmp[5201]*kernel[7]+tmp[5202]*kernel[8];
				ans[5102]<=tmp[5001]*kernel[0]+tmp[5002]*kernel[1]+tmp[5003]*kernel[2]+tmp[5101]*kernel[3]+tmp[5102]*kernel[4]+tmp[5103]*kernel[5]+tmp[5201]*kernel[6]+tmp[5202]*kernel[7]+tmp[5203]*kernel[8];
				ans[5103]<=tmp[5002]*kernel[0]+tmp[5003]*kernel[1]+tmp[5004]*kernel[2]+tmp[5102]*kernel[3]+tmp[5103]*kernel[4]+tmp[5104]*kernel[5]+tmp[5202]*kernel[6]+tmp[5203]*kernel[7]+tmp[5204]*kernel[8];
				ans[5104]<=tmp[5003]*kernel[0]+tmp[5004]*kernel[1]+tmp[5005]*kernel[2]+tmp[5103]*kernel[3]+tmp[5104]*kernel[4]+tmp[5105]*kernel[5]+tmp[5203]*kernel[6]+tmp[5204]*kernel[7]+tmp[5205]*kernel[8];
				ans[5105]<=tmp[5004]*kernel[0]+tmp[5005]*kernel[1]+tmp[5006]*kernel[2]+tmp[5104]*kernel[3]+tmp[5105]*kernel[4]+tmp[5106]*kernel[5]+tmp[5204]*kernel[6]+tmp[5205]*kernel[7]+tmp[5206]*kernel[8];
				ans[5106]<=tmp[5005]*kernel[0]+tmp[5006]*kernel[1]+tmp[5007]*kernel[2]+tmp[5105]*kernel[3]+tmp[5106]*kernel[4]+tmp[5107]*kernel[5]+tmp[5205]*kernel[6]+tmp[5206]*kernel[7]+tmp[5207]*kernel[8];
				ans[5107]<=tmp[5006]*kernel[0]+tmp[5007]*kernel[1]+tmp[5008]*kernel[2]+tmp[5106]*kernel[3]+tmp[5107]*kernel[4]+tmp[5108]*kernel[5]+tmp[5206]*kernel[6]+tmp[5207]*kernel[7]+tmp[5208]*kernel[8];
				ans[5108]<=tmp[5007]*kernel[0]+tmp[5008]*kernel[1]+tmp[5009]*kernel[2]+tmp[5107]*kernel[3]+tmp[5108]*kernel[4]+tmp[5109]*kernel[5]+tmp[5207]*kernel[6]+tmp[5208]*kernel[7]+tmp[5209]*kernel[8];
				ans[5109]<=tmp[5008]*kernel[0]+tmp[5009]*kernel[1]+tmp[5010]*kernel[2]+tmp[5108]*kernel[3]+tmp[5109]*kernel[4]+tmp[5110]*kernel[5]+tmp[5208]*kernel[6]+tmp[5209]*kernel[7]+tmp[5210]*kernel[8];
				ans[5110]<=tmp[5009]*kernel[0]+tmp[5010]*kernel[1]+tmp[5011]*kernel[2]+tmp[5109]*kernel[3]+tmp[5110]*kernel[4]+tmp[5111]*kernel[5]+tmp[5209]*kernel[6]+tmp[5210]*kernel[7]+tmp[5211]*kernel[8];
				ans[5111]<=tmp[5010]*kernel[0]+tmp[5011]*kernel[1]+tmp[5012]*kernel[2]+tmp[5110]*kernel[3]+tmp[5111]*kernel[4]+tmp[5112]*kernel[5]+tmp[5210]*kernel[6]+tmp[5211]*kernel[7]+tmp[5212]*kernel[8];
				ans[5112]<=tmp[5011]*kernel[0]+tmp[5012]*kernel[1]+tmp[5013]*kernel[2]+tmp[5111]*kernel[3]+tmp[5112]*kernel[4]+tmp[5113]*kernel[5]+tmp[5211]*kernel[6]+tmp[5212]*kernel[7]+tmp[5213]*kernel[8];
				ans[5113]<=tmp[5012]*kernel[0]+tmp[5013]*kernel[1]+tmp[5014]*kernel[2]+tmp[5112]*kernel[3]+tmp[5113]*kernel[4]+tmp[5114]*kernel[5]+tmp[5212]*kernel[6]+tmp[5213]*kernel[7]+tmp[5214]*kernel[8];
				ans[5114]<=tmp[5013]*kernel[0]+tmp[5014]*kernel[1]+tmp[5015]*kernel[2]+tmp[5113]*kernel[3]+tmp[5114]*kernel[4]+tmp[5115]*kernel[5]+tmp[5213]*kernel[6]+tmp[5214]*kernel[7]+tmp[5215]*kernel[8];
				ans[5115]<=tmp[5014]*kernel[0]+tmp[5015]*kernel[1]+tmp[5016]*kernel[2]+tmp[5114]*kernel[3]+tmp[5115]*kernel[4]+tmp[5116]*kernel[5]+tmp[5214]*kernel[6]+tmp[5215]*kernel[7]+tmp[5216]*kernel[8];
				ans[5116]<=tmp[5015]*kernel[0]+tmp[5016]*kernel[1]+tmp[5017]*kernel[2]+tmp[5115]*kernel[3]+tmp[5116]*kernel[4]+tmp[5117]*kernel[5]+tmp[5215]*kernel[6]+tmp[5216]*kernel[7]+tmp[5217]*kernel[8];
				ans[5117]<=tmp[5016]*kernel[0]+tmp[5017]*kernel[1]+tmp[5018]*kernel[2]+tmp[5116]*kernel[3]+tmp[5117]*kernel[4]+tmp[5118]*kernel[5]+tmp[5216]*kernel[6]+tmp[5217]*kernel[7]+tmp[5218]*kernel[8];
				ans[5118]<=tmp[5017]*kernel[0]+tmp[5018]*kernel[1]+tmp[5019]*kernel[2]+tmp[5117]*kernel[3]+tmp[5118]*kernel[4]+tmp[5119]*kernel[5]+tmp[5217]*kernel[6]+tmp[5218]*kernel[7]+tmp[5219]*kernel[8];
				ans[5119]<=tmp[5018]*kernel[0]+tmp[5019]*kernel[1]+tmp[5020]*kernel[2]+tmp[5118]*kernel[3]+tmp[5119]*kernel[4]+tmp[5120]*kernel[5]+tmp[5218]*kernel[6]+tmp[5219]*kernel[7]+tmp[5220]*kernel[8];
				ans[5120]<=tmp[5019]*kernel[0]+tmp[5020]*kernel[1]+tmp[5021]*kernel[2]+tmp[5119]*kernel[3]+tmp[5120]*kernel[4]+tmp[5121]*kernel[5]+tmp[5219]*kernel[6]+tmp[5220]*kernel[7]+tmp[5221]*kernel[8];
				ans[5121]<=tmp[5020]*kernel[0]+tmp[5021]*kernel[1]+tmp[5022]*kernel[2]+tmp[5120]*kernel[3]+tmp[5121]*kernel[4]+tmp[5122]*kernel[5]+tmp[5220]*kernel[6]+tmp[5221]*kernel[7]+tmp[5222]*kernel[8];
				ans[5122]<=tmp[5021]*kernel[0]+tmp[5022]*kernel[1]+tmp[5023]*kernel[2]+tmp[5121]*kernel[3]+tmp[5122]*kernel[4]+tmp[5123]*kernel[5]+tmp[5221]*kernel[6]+tmp[5222]*kernel[7]+tmp[5223]*kernel[8];
				ans[5123]<=tmp[5022]*kernel[0]+tmp[5023]*kernel[1]+tmp[5024]*kernel[2]+tmp[5122]*kernel[3]+tmp[5123]*kernel[4]+tmp[5124]*kernel[5]+tmp[5222]*kernel[6]+tmp[5223]*kernel[7]+tmp[5224]*kernel[8];
				ans[5124]<=tmp[5023]*kernel[0]+tmp[5024]*kernel[1]+tmp[5025]*kernel[2]+tmp[5123]*kernel[3]+tmp[5124]*kernel[4]+tmp[5125]*kernel[5]+tmp[5223]*kernel[6]+tmp[5224]*kernel[7]+tmp[5225]*kernel[8];
				ans[5125]<=tmp[5024]*kernel[0]+tmp[5025]*kernel[1]+tmp[5026]*kernel[2]+tmp[5124]*kernel[3]+tmp[5125]*kernel[4]+tmp[5126]*kernel[5]+tmp[5224]*kernel[6]+tmp[5225]*kernel[7]+tmp[5226]*kernel[8];
				ans[5126]<=tmp[5025]*kernel[0]+tmp[5026]*kernel[1]+tmp[5027]*kernel[2]+tmp[5125]*kernel[3]+tmp[5126]*kernel[4]+tmp[5127]*kernel[5]+tmp[5225]*kernel[6]+tmp[5226]*kernel[7]+tmp[5227]*kernel[8];
				ans[5127]<=tmp[5026]*kernel[0]+tmp[5027]*kernel[1]+tmp[5028]*kernel[2]+tmp[5126]*kernel[3]+tmp[5127]*kernel[4]+tmp[5128]*kernel[5]+tmp[5226]*kernel[6]+tmp[5227]*kernel[7]+tmp[5228]*kernel[8];
				ans[5128]<=tmp[5027]*kernel[0]+tmp[5028]*kernel[1]+tmp[5029]*kernel[2]+tmp[5127]*kernel[3]+tmp[5128]*kernel[4]+tmp[5129]*kernel[5]+tmp[5227]*kernel[6]+tmp[5228]*kernel[7]+tmp[5229]*kernel[8];
				ans[5129]<=tmp[5028]*kernel[0]+tmp[5029]*kernel[1]+tmp[5030]*kernel[2]+tmp[5128]*kernel[3]+tmp[5129]*kernel[4]+tmp[5130]*kernel[5]+tmp[5228]*kernel[6]+tmp[5229]*kernel[7]+tmp[5230]*kernel[8];
				ans[5130]<=tmp[5029]*kernel[0]+tmp[5030]*kernel[1]+tmp[5031]*kernel[2]+tmp[5129]*kernel[3]+tmp[5130]*kernel[4]+tmp[5131]*kernel[5]+tmp[5229]*kernel[6]+tmp[5230]*kernel[7]+tmp[5231]*kernel[8];
				ans[5131]<=tmp[5030]*kernel[0]+tmp[5031]*kernel[1]+tmp[5032]*kernel[2]+tmp[5130]*kernel[3]+tmp[5131]*kernel[4]+tmp[5132]*kernel[5]+tmp[5230]*kernel[6]+tmp[5231]*kernel[7]+tmp[5232]*kernel[8];
				ans[5132]<=tmp[5031]*kernel[0]+tmp[5032]*kernel[1]+tmp[5033]*kernel[2]+tmp[5131]*kernel[3]+tmp[5132]*kernel[4]+tmp[5133]*kernel[5]+tmp[5231]*kernel[6]+tmp[5232]*kernel[7]+tmp[5233]*kernel[8];
				ans[5133]<=tmp[5032]*kernel[0]+tmp[5033]*kernel[1]+tmp[5034]*kernel[2]+tmp[5132]*kernel[3]+tmp[5133]*kernel[4]+tmp[5134]*kernel[5]+tmp[5232]*kernel[6]+tmp[5233]*kernel[7]+tmp[5234]*kernel[8];
				ans[5134]<=tmp[5033]*kernel[0]+tmp[5034]*kernel[1]+tmp[5035]*kernel[2]+tmp[5133]*kernel[3]+tmp[5134]*kernel[4]+tmp[5135]*kernel[5]+tmp[5233]*kernel[6]+tmp[5234]*kernel[7]+tmp[5235]*kernel[8];
				ans[5135]<=tmp[5034]*kernel[0]+tmp[5035]*kernel[1]+tmp[5036]*kernel[2]+tmp[5134]*kernel[3]+tmp[5135]*kernel[4]+tmp[5136]*kernel[5]+tmp[5234]*kernel[6]+tmp[5235]*kernel[7]+tmp[5236]*kernel[8];
				ans[5136]<=tmp[5035]*kernel[0]+tmp[5036]*kernel[1]+tmp[5037]*kernel[2]+tmp[5135]*kernel[3]+tmp[5136]*kernel[4]+tmp[5137]*kernel[5]+tmp[5235]*kernel[6]+tmp[5236]*kernel[7]+tmp[5237]*kernel[8];
				ans[5137]<=tmp[5036]*kernel[0]+tmp[5037]*kernel[1]+tmp[5038]*kernel[2]+tmp[5136]*kernel[3]+tmp[5137]*kernel[4]+tmp[5138]*kernel[5]+tmp[5236]*kernel[6]+tmp[5237]*kernel[7]+tmp[5238]*kernel[8];
				ans[5138]<=tmp[5037]*kernel[0]+tmp[5038]*kernel[1]+tmp[5039]*kernel[2]+tmp[5137]*kernel[3]+tmp[5138]*kernel[4]+tmp[5139]*kernel[5]+tmp[5237]*kernel[6]+tmp[5238]*kernel[7]+tmp[5239]*kernel[8];
				ans[5139]<=tmp[5038]*kernel[0]+tmp[5039]*kernel[1]+tmp[5040]*kernel[2]+tmp[5138]*kernel[3]+tmp[5139]*kernel[4]+tmp[5140]*kernel[5]+tmp[5238]*kernel[6]+tmp[5239]*kernel[7]+tmp[5240]*kernel[8];
				ans[5140]<=tmp[5039]*kernel[0]+tmp[5040]*kernel[1]+tmp[5041]*kernel[2]+tmp[5139]*kernel[3]+tmp[5140]*kernel[4]+tmp[5141]*kernel[5]+tmp[5239]*kernel[6]+tmp[5240]*kernel[7]+tmp[5241]*kernel[8];
				ans[5141]<=tmp[5040]*kernel[0]+tmp[5041]*kernel[1]+tmp[5042]*kernel[2]+tmp[5140]*kernel[3]+tmp[5141]*kernel[4]+tmp[5142]*kernel[5]+tmp[5240]*kernel[6]+tmp[5241]*kernel[7]+tmp[5242]*kernel[8];
				ans[5142]<=tmp[5041]*kernel[0]+tmp[5042]*kernel[1]+tmp[5043]*kernel[2]+tmp[5141]*kernel[3]+tmp[5142]*kernel[4]+tmp[5143]*kernel[5]+tmp[5241]*kernel[6]+tmp[5242]*kernel[7]+tmp[5243]*kernel[8];
				ans[5143]<=tmp[5042]*kernel[0]+tmp[5043]*kernel[1]+tmp[5044]*kernel[2]+tmp[5142]*kernel[3]+tmp[5143]*kernel[4]+tmp[5144]*kernel[5]+tmp[5242]*kernel[6]+tmp[5243]*kernel[7]+tmp[5244]*kernel[8];
				ans[5144]<=tmp[5043]*kernel[0]+tmp[5044]*kernel[1]+tmp[5045]*kernel[2]+tmp[5143]*kernel[3]+tmp[5144]*kernel[4]+tmp[5145]*kernel[5]+tmp[5243]*kernel[6]+tmp[5244]*kernel[7]+tmp[5245]*kernel[8];
				ans[5145]<=tmp[5044]*kernel[0]+tmp[5045]*kernel[1]+tmp[5046]*kernel[2]+tmp[5144]*kernel[3]+tmp[5145]*kernel[4]+tmp[5146]*kernel[5]+tmp[5244]*kernel[6]+tmp[5245]*kernel[7]+tmp[5246]*kernel[8];
				ans[5146]<=tmp[5045]*kernel[0]+tmp[5046]*kernel[1]+tmp[5047]*kernel[2]+tmp[5145]*kernel[3]+tmp[5146]*kernel[4]+tmp[5147]*kernel[5]+tmp[5245]*kernel[6]+tmp[5246]*kernel[7]+tmp[5247]*kernel[8];
				ans[5147]<=tmp[5046]*kernel[0]+tmp[5047]*kernel[1]+tmp[5048]*kernel[2]+tmp[5146]*kernel[3]+tmp[5147]*kernel[4]+tmp[5148]*kernel[5]+tmp[5246]*kernel[6]+tmp[5247]*kernel[7]+tmp[5248]*kernel[8];
				ans[5148]<=tmp[5047]*kernel[0]+tmp[5048]*kernel[1]+tmp[5049]*kernel[2]+tmp[5147]*kernel[3]+tmp[5148]*kernel[4]+tmp[5149]*kernel[5]+tmp[5247]*kernel[6]+tmp[5248]*kernel[7]+tmp[5249]*kernel[8];
				ans[5149]<=tmp[5048]*kernel[0]+tmp[5049]*kernel[1]+tmp[5050]*kernel[2]+tmp[5148]*kernel[3]+tmp[5149]*kernel[4]+tmp[5150]*kernel[5]+tmp[5248]*kernel[6]+tmp[5249]*kernel[7]+tmp[5250]*kernel[8];
				ans[5150]<=tmp[5049]*kernel[0]+tmp[5050]*kernel[1]+tmp[5051]*kernel[2]+tmp[5149]*kernel[3]+tmp[5150]*kernel[4]+tmp[5151]*kernel[5]+tmp[5249]*kernel[6]+tmp[5250]*kernel[7]+tmp[5251]*kernel[8];
				ans[5151]<=tmp[5050]*kernel[0]+tmp[5051]*kernel[1]+tmp[5052]*kernel[2]+tmp[5150]*kernel[3]+tmp[5151]*kernel[4]+tmp[5152]*kernel[5]+tmp[5250]*kernel[6]+tmp[5251]*kernel[7]+tmp[5252]*kernel[8];
				ans[5152]<=tmp[5051]*kernel[0]+tmp[5052]*kernel[1]+tmp[5053]*kernel[2]+tmp[5151]*kernel[3]+tmp[5152]*kernel[4]+tmp[5153]*kernel[5]+tmp[5251]*kernel[6]+tmp[5252]*kernel[7]+tmp[5253]*kernel[8];
				ans[5153]<=tmp[5052]*kernel[0]+tmp[5053]*kernel[1]+tmp[5054]*kernel[2]+tmp[5152]*kernel[3]+tmp[5153]*kernel[4]+tmp[5154]*kernel[5]+tmp[5252]*kernel[6]+tmp[5253]*kernel[7]+tmp[5254]*kernel[8];
				ans[5154]<=tmp[5053]*kernel[0]+tmp[5054]*kernel[1]+tmp[5055]*kernel[2]+tmp[5153]*kernel[3]+tmp[5154]*kernel[4]+tmp[5155]*kernel[5]+tmp[5253]*kernel[6]+tmp[5254]*kernel[7]+tmp[5255]*kernel[8];
				ans[5155]<=tmp[5054]*kernel[0]+tmp[5055]*kernel[1]+tmp[5056]*kernel[2]+tmp[5154]*kernel[3]+tmp[5155]*kernel[4]+tmp[5156]*kernel[5]+tmp[5254]*kernel[6]+tmp[5255]*kernel[7]+tmp[5256]*kernel[8];
				ans[5156]<=tmp[5055]*kernel[0]+tmp[5056]*kernel[1]+tmp[5057]*kernel[2]+tmp[5155]*kernel[3]+tmp[5156]*kernel[4]+tmp[5157]*kernel[5]+tmp[5255]*kernel[6]+tmp[5256]*kernel[7]+tmp[5257]*kernel[8];
				ans[5157]<=tmp[5056]*kernel[0]+tmp[5057]*kernel[1]+tmp[5058]*kernel[2]+tmp[5156]*kernel[3]+tmp[5157]*kernel[4]+tmp[5158]*kernel[5]+tmp[5256]*kernel[6]+tmp[5257]*kernel[7]+tmp[5258]*kernel[8];
				ans[5158]<=tmp[5057]*kernel[0]+tmp[5058]*kernel[1]+tmp[5059]*kernel[2]+tmp[5157]*kernel[3]+tmp[5158]*kernel[4]+tmp[5159]*kernel[5]+tmp[5257]*kernel[6]+tmp[5258]*kernel[7]+tmp[5259]*kernel[8];
				ans[5159]<=tmp[5058]*kernel[0]+tmp[5059]*kernel[1]+tmp[5060]*kernel[2]+tmp[5158]*kernel[3]+tmp[5159]*kernel[4]+tmp[5160]*kernel[5]+tmp[5258]*kernel[6]+tmp[5259]*kernel[7]+tmp[5260]*kernel[8];
				ans[5160]<=tmp[5059]*kernel[0]+tmp[5060]*kernel[1]+tmp[5061]*kernel[2]+tmp[5159]*kernel[3]+tmp[5160]*kernel[4]+tmp[5161]*kernel[5]+tmp[5259]*kernel[6]+tmp[5260]*kernel[7]+tmp[5261]*kernel[8];
				ans[5161]<=tmp[5060]*kernel[0]+tmp[5061]*kernel[1]+tmp[5062]*kernel[2]+tmp[5160]*kernel[3]+tmp[5161]*kernel[4]+tmp[5162]*kernel[5]+tmp[5260]*kernel[6]+tmp[5261]*kernel[7]+tmp[5262]*kernel[8];
				ans[5162]<=tmp[5061]*kernel[0]+tmp[5062]*kernel[1]+tmp[5063]*kernel[2]+tmp[5161]*kernel[3]+tmp[5162]*kernel[4]+tmp[5163]*kernel[5]+tmp[5261]*kernel[6]+tmp[5262]*kernel[7]+tmp[5263]*kernel[8];
				ans[5163]<=tmp[5062]*kernel[0]+tmp[5063]*kernel[1]+tmp[5064]*kernel[2]+tmp[5162]*kernel[3]+tmp[5163]*kernel[4]+tmp[5164]*kernel[5]+tmp[5262]*kernel[6]+tmp[5263]*kernel[7]+tmp[5264]*kernel[8];
				ans[5164]<=tmp[5063]*kernel[0]+tmp[5064]*kernel[1]+tmp[5065]*kernel[2]+tmp[5163]*kernel[3]+tmp[5164]*kernel[4]+tmp[5165]*kernel[5]+tmp[5263]*kernel[6]+tmp[5264]*kernel[7]+tmp[5265]*kernel[8];
				ans[5165]<=tmp[5064]*kernel[0]+tmp[5065]*kernel[1]+tmp[5066]*kernel[2]+tmp[5164]*kernel[3]+tmp[5165]*kernel[4]+tmp[5166]*kernel[5]+tmp[5264]*kernel[6]+tmp[5265]*kernel[7]+tmp[5266]*kernel[8];
				ans[5166]<=tmp[5065]*kernel[0]+tmp[5066]*kernel[1]+tmp[5067]*kernel[2]+tmp[5165]*kernel[3]+tmp[5166]*kernel[4]+tmp[5167]*kernel[5]+tmp[5265]*kernel[6]+tmp[5266]*kernel[7]+tmp[5267]*kernel[8];
				ans[5167]<=tmp[5066]*kernel[0]+tmp[5067]*kernel[1]+tmp[5068]*kernel[2]+tmp[5166]*kernel[3]+tmp[5167]*kernel[4]+tmp[5168]*kernel[5]+tmp[5266]*kernel[6]+tmp[5267]*kernel[7]+tmp[5268]*kernel[8];
				ans[5168]<=tmp[5067]*kernel[0]+tmp[5068]*kernel[1]+tmp[5069]*kernel[2]+tmp[5167]*kernel[3]+tmp[5168]*kernel[4]+tmp[5169]*kernel[5]+tmp[5267]*kernel[6]+tmp[5268]*kernel[7]+tmp[5269]*kernel[8];
				ans[5169]<=tmp[5068]*kernel[0]+tmp[5069]*kernel[1]+tmp[5070]*kernel[2]+tmp[5168]*kernel[3]+tmp[5169]*kernel[4]+tmp[5170]*kernel[5]+tmp[5268]*kernel[6]+tmp[5269]*kernel[7]+tmp[5270]*kernel[8];
				ans[5170]<=tmp[5069]*kernel[0]+tmp[5070]*kernel[1]+tmp[5071]*kernel[2]+tmp[5169]*kernel[3]+tmp[5170]*kernel[4]+tmp[5171]*kernel[5]+tmp[5269]*kernel[6]+tmp[5270]*kernel[7]+tmp[5271]*kernel[8];
				ans[5171]<=tmp[5070]*kernel[0]+tmp[5071]*kernel[1]+tmp[5072]*kernel[2]+tmp[5170]*kernel[3]+tmp[5171]*kernel[4]+tmp[5172]*kernel[5]+tmp[5270]*kernel[6]+tmp[5271]*kernel[7]+tmp[5272]*kernel[8];
				ans[5172]<=tmp[5071]*kernel[0]+tmp[5072]*kernel[1]+tmp[5073]*kernel[2]+tmp[5171]*kernel[3]+tmp[5172]*kernel[4]+tmp[5173]*kernel[5]+tmp[5271]*kernel[6]+tmp[5272]*kernel[7]+tmp[5273]*kernel[8];
				ans[5173]<=tmp[5072]*kernel[0]+tmp[5073]*kernel[1]+tmp[5074]*kernel[2]+tmp[5172]*kernel[3]+tmp[5173]*kernel[4]+tmp[5174]*kernel[5]+tmp[5272]*kernel[6]+tmp[5273]*kernel[7]+tmp[5274]*kernel[8];
				ans[5174]<=tmp[5073]*kernel[0]+tmp[5074]*kernel[1]+tmp[5075]*kernel[2]+tmp[5173]*kernel[3]+tmp[5174]*kernel[4]+tmp[5175]*kernel[5]+tmp[5273]*kernel[6]+tmp[5274]*kernel[7]+tmp[5275]*kernel[8];
				ans[5175]<=tmp[5074]*kernel[0]+tmp[5075]*kernel[1]+tmp[5076]*kernel[2]+tmp[5174]*kernel[3]+tmp[5175]*kernel[4]+tmp[5176]*kernel[5]+tmp[5274]*kernel[6]+tmp[5275]*kernel[7]+tmp[5276]*kernel[8];
				ans[5176]<=tmp[5075]*kernel[0]+tmp[5076]*kernel[1]+tmp[5077]*kernel[2]+tmp[5175]*kernel[3]+tmp[5176]*kernel[4]+tmp[5177]*kernel[5]+tmp[5275]*kernel[6]+tmp[5276]*kernel[7]+tmp[5277]*kernel[8];
				ans[5177]<=tmp[5076]*kernel[0]+tmp[5077]*kernel[1]+tmp[5078]*kernel[2]+tmp[5176]*kernel[3]+tmp[5177]*kernel[4]+tmp[5178]*kernel[5]+tmp[5276]*kernel[6]+tmp[5277]*kernel[7]+tmp[5278]*kernel[8];
				ans[5178]<=tmp[5077]*kernel[0]+tmp[5078]*kernel[1]+tmp[5079]*kernel[2]+tmp[5177]*kernel[3]+tmp[5178]*kernel[4]+tmp[5179]*kernel[5]+tmp[5277]*kernel[6]+tmp[5278]*kernel[7]+tmp[5279]*kernel[8];
				ans[5179]<=tmp[5078]*kernel[0]+tmp[5079]*kernel[1]+tmp[5080]*kernel[2]+tmp[5178]*kernel[3]+tmp[5179]*kernel[4]+tmp[5180]*kernel[5]+tmp[5278]*kernel[6]+tmp[5279]*kernel[7]+tmp[5280]*kernel[8];
				ans[5180]<=tmp[5079]*kernel[0]+tmp[5080]*kernel[1]+tmp[5081]*kernel[2]+tmp[5179]*kernel[3]+tmp[5180]*kernel[4]+tmp[5181]*kernel[5]+tmp[5279]*kernel[6]+tmp[5280]*kernel[7]+tmp[5281]*kernel[8];
				ans[5181]<=tmp[5080]*kernel[0]+tmp[5081]*kernel[1]+tmp[5082]*kernel[2]+tmp[5180]*kernel[3]+tmp[5181]*kernel[4]+tmp[5182]*kernel[5]+tmp[5280]*kernel[6]+tmp[5281]*kernel[7]+tmp[5282]*kernel[8];
				ans[5182]<=tmp[5081]*kernel[0]+tmp[5082]*kernel[1]+tmp[5083]*kernel[2]+tmp[5181]*kernel[3]+tmp[5182]*kernel[4]+tmp[5183]*kernel[5]+tmp[5281]*kernel[6]+tmp[5282]*kernel[7]+tmp[5283]*kernel[8];
				ans[5183]<=tmp[5082]*kernel[0]+tmp[5083]*kernel[1]+tmp[5084]*kernel[2]+tmp[5182]*kernel[3]+tmp[5183]*kernel[4]+tmp[5184]*kernel[5]+tmp[5282]*kernel[6]+tmp[5283]*kernel[7]+tmp[5284]*kernel[8];
				ans[5184]<=tmp[5083]*kernel[0]+tmp[5084]*kernel[1]+tmp[5085]*kernel[2]+tmp[5183]*kernel[3]+tmp[5184]*kernel[4]+tmp[5185]*kernel[5]+tmp[5283]*kernel[6]+tmp[5284]*kernel[7]+tmp[5285]*kernel[8];
				ans[5185]<=tmp[5084]*kernel[0]+tmp[5085]*kernel[1]+tmp[5086]*kernel[2]+tmp[5184]*kernel[3]+tmp[5185]*kernel[4]+tmp[5186]*kernel[5]+tmp[5284]*kernel[6]+tmp[5285]*kernel[7]+tmp[5286]*kernel[8];
				ans[5186]<=tmp[5085]*kernel[0]+tmp[5086]*kernel[1]+tmp[5087]*kernel[2]+tmp[5185]*kernel[3]+tmp[5186]*kernel[4]+tmp[5187]*kernel[5]+tmp[5285]*kernel[6]+tmp[5286]*kernel[7]+tmp[5287]*kernel[8];
				ans[5187]<=tmp[5086]*kernel[0]+tmp[5087]*kernel[1]+tmp[5088]*kernel[2]+tmp[5186]*kernel[3]+tmp[5187]*kernel[4]+tmp[5188]*kernel[5]+tmp[5286]*kernel[6]+tmp[5287]*kernel[7]+tmp[5288]*kernel[8];
				ans[5188]<=tmp[5087]*kernel[0]+tmp[5088]*kernel[1]+tmp[5089]*kernel[2]+tmp[5187]*kernel[3]+tmp[5188]*kernel[4]+tmp[5189]*kernel[5]+tmp[5287]*kernel[6]+tmp[5288]*kernel[7]+tmp[5289]*kernel[8];
				ans[5189]<=tmp[5088]*kernel[0]+tmp[5089]*kernel[1]+tmp[5090]*kernel[2]+tmp[5188]*kernel[3]+tmp[5189]*kernel[4]+tmp[5190]*kernel[5]+tmp[5288]*kernel[6]+tmp[5289]*kernel[7]+tmp[5290]*kernel[8];
				ans[5190]<=tmp[5089]*kernel[0]+tmp[5090]*kernel[1]+tmp[5091]*kernel[2]+tmp[5189]*kernel[3]+tmp[5190]*kernel[4]+tmp[5191]*kernel[5]+tmp[5289]*kernel[6]+tmp[5290]*kernel[7]+tmp[5291]*kernel[8];
				ans[5191]<=tmp[5090]*kernel[0]+tmp[5091]*kernel[1]+tmp[5092]*kernel[2]+tmp[5190]*kernel[3]+tmp[5191]*kernel[4]+tmp[5192]*kernel[5]+tmp[5290]*kernel[6]+tmp[5291]*kernel[7]+tmp[5292]*kernel[8];
				ans[5192]<=tmp[5091]*kernel[0]+tmp[5092]*kernel[1]+tmp[5093]*kernel[2]+tmp[5191]*kernel[3]+tmp[5192]*kernel[4]+tmp[5193]*kernel[5]+tmp[5291]*kernel[6]+tmp[5292]*kernel[7]+tmp[5293]*kernel[8];
				ans[5193]<=tmp[5092]*kernel[0]+tmp[5093]*kernel[1]+tmp[5094]*kernel[2]+tmp[5192]*kernel[3]+tmp[5193]*kernel[4]+tmp[5194]*kernel[5]+tmp[5292]*kernel[6]+tmp[5293]*kernel[7]+tmp[5294]*kernel[8];
				ans[5194]<=tmp[5093]*kernel[0]+tmp[5094]*kernel[1]+tmp[5095]*kernel[2]+tmp[5193]*kernel[3]+tmp[5194]*kernel[4]+tmp[5195]*kernel[5]+tmp[5293]*kernel[6]+tmp[5294]*kernel[7]+tmp[5295]*kernel[8];
				ans[5195]<=tmp[5094]*kernel[0]+tmp[5095]*kernel[1]+tmp[5096]*kernel[2]+tmp[5194]*kernel[3]+tmp[5195]*kernel[4]+tmp[5196]*kernel[5]+tmp[5294]*kernel[6]+tmp[5295]*kernel[7]+tmp[5296]*kernel[8];
				ans[5196]<=tmp[5095]*kernel[0]+tmp[5096]*kernel[1]+tmp[5097]*kernel[2]+tmp[5195]*kernel[3]+tmp[5196]*kernel[4]+tmp[5197]*kernel[5]+tmp[5295]*kernel[6]+tmp[5296]*kernel[7]+tmp[5297]*kernel[8];
				ans[5197]<=tmp[5096]*kernel[0]+tmp[5097]*kernel[1]+tmp[5098]*kernel[2]+tmp[5196]*kernel[3]+tmp[5197]*kernel[4]+tmp[5198]*kernel[5]+tmp[5296]*kernel[6]+tmp[5297]*kernel[7]+tmp[5298]*kernel[8];
				ans[5198]<=tmp[5097]*kernel[0]+tmp[5098]*kernel[1]+tmp[5099]*kernel[2]+tmp[5197]*kernel[3]+tmp[5198]*kernel[4]+tmp[5199]*kernel[5]+tmp[5297]*kernel[6]+tmp[5298]*kernel[7]+tmp[5299]*kernel[8];
				ans[5199]<=tmp[5098]*kernel[0]+tmp[5099]*kernel[1]+tmp[5198]*kernel[3]+tmp[5199]*kernel[4]+tmp[5298]*kernel[6]+tmp[5299]*kernel[7];
				ans[5200]<=tmp[5100]*kernel[1]+tmp[5101]*kernel[2]+tmp[5200]*kernel[4]+tmp[5201]*kernel[5]+tmp[5300]*kernel[7]+tmp[5301]*kernel[8];
				ans[5201]<=tmp[5100]*kernel[0]+tmp[5101]*kernel[1]+tmp[5102]*kernel[2]+tmp[5200]*kernel[3]+tmp[5201]*kernel[4]+tmp[5202]*kernel[5]+tmp[5300]*kernel[6]+tmp[5301]*kernel[7]+tmp[5302]*kernel[8];
				ans[5202]<=tmp[5101]*kernel[0]+tmp[5102]*kernel[1]+tmp[5103]*kernel[2]+tmp[5201]*kernel[3]+tmp[5202]*kernel[4]+tmp[5203]*kernel[5]+tmp[5301]*kernel[6]+tmp[5302]*kernel[7]+tmp[5303]*kernel[8];
				ans[5203]<=tmp[5102]*kernel[0]+tmp[5103]*kernel[1]+tmp[5104]*kernel[2]+tmp[5202]*kernel[3]+tmp[5203]*kernel[4]+tmp[5204]*kernel[5]+tmp[5302]*kernel[6]+tmp[5303]*kernel[7]+tmp[5304]*kernel[8];
				ans[5204]<=tmp[5103]*kernel[0]+tmp[5104]*kernel[1]+tmp[5105]*kernel[2]+tmp[5203]*kernel[3]+tmp[5204]*kernel[4]+tmp[5205]*kernel[5]+tmp[5303]*kernel[6]+tmp[5304]*kernel[7]+tmp[5305]*kernel[8];
				ans[5205]<=tmp[5104]*kernel[0]+tmp[5105]*kernel[1]+tmp[5106]*kernel[2]+tmp[5204]*kernel[3]+tmp[5205]*kernel[4]+tmp[5206]*kernel[5]+tmp[5304]*kernel[6]+tmp[5305]*kernel[7]+tmp[5306]*kernel[8];
				ans[5206]<=tmp[5105]*kernel[0]+tmp[5106]*kernel[1]+tmp[5107]*kernel[2]+tmp[5205]*kernel[3]+tmp[5206]*kernel[4]+tmp[5207]*kernel[5]+tmp[5305]*kernel[6]+tmp[5306]*kernel[7]+tmp[5307]*kernel[8];
				ans[5207]<=tmp[5106]*kernel[0]+tmp[5107]*kernel[1]+tmp[5108]*kernel[2]+tmp[5206]*kernel[3]+tmp[5207]*kernel[4]+tmp[5208]*kernel[5]+tmp[5306]*kernel[6]+tmp[5307]*kernel[7]+tmp[5308]*kernel[8];
				ans[5208]<=tmp[5107]*kernel[0]+tmp[5108]*kernel[1]+tmp[5109]*kernel[2]+tmp[5207]*kernel[3]+tmp[5208]*kernel[4]+tmp[5209]*kernel[5]+tmp[5307]*kernel[6]+tmp[5308]*kernel[7]+tmp[5309]*kernel[8];
				ans[5209]<=tmp[5108]*kernel[0]+tmp[5109]*kernel[1]+tmp[5110]*kernel[2]+tmp[5208]*kernel[3]+tmp[5209]*kernel[4]+tmp[5210]*kernel[5]+tmp[5308]*kernel[6]+tmp[5309]*kernel[7]+tmp[5310]*kernel[8];
				ans[5210]<=tmp[5109]*kernel[0]+tmp[5110]*kernel[1]+tmp[5111]*kernel[2]+tmp[5209]*kernel[3]+tmp[5210]*kernel[4]+tmp[5211]*kernel[5]+tmp[5309]*kernel[6]+tmp[5310]*kernel[7]+tmp[5311]*kernel[8];
				ans[5211]<=tmp[5110]*kernel[0]+tmp[5111]*kernel[1]+tmp[5112]*kernel[2]+tmp[5210]*kernel[3]+tmp[5211]*kernel[4]+tmp[5212]*kernel[5]+tmp[5310]*kernel[6]+tmp[5311]*kernel[7]+tmp[5312]*kernel[8];
				ans[5212]<=tmp[5111]*kernel[0]+tmp[5112]*kernel[1]+tmp[5113]*kernel[2]+tmp[5211]*kernel[3]+tmp[5212]*kernel[4]+tmp[5213]*kernel[5]+tmp[5311]*kernel[6]+tmp[5312]*kernel[7]+tmp[5313]*kernel[8];
				ans[5213]<=tmp[5112]*kernel[0]+tmp[5113]*kernel[1]+tmp[5114]*kernel[2]+tmp[5212]*kernel[3]+tmp[5213]*kernel[4]+tmp[5214]*kernel[5]+tmp[5312]*kernel[6]+tmp[5313]*kernel[7]+tmp[5314]*kernel[8];
				ans[5214]<=tmp[5113]*kernel[0]+tmp[5114]*kernel[1]+tmp[5115]*kernel[2]+tmp[5213]*kernel[3]+tmp[5214]*kernel[4]+tmp[5215]*kernel[5]+tmp[5313]*kernel[6]+tmp[5314]*kernel[7]+tmp[5315]*kernel[8];
				ans[5215]<=tmp[5114]*kernel[0]+tmp[5115]*kernel[1]+tmp[5116]*kernel[2]+tmp[5214]*kernel[3]+tmp[5215]*kernel[4]+tmp[5216]*kernel[5]+tmp[5314]*kernel[6]+tmp[5315]*kernel[7]+tmp[5316]*kernel[8];
				ans[5216]<=tmp[5115]*kernel[0]+tmp[5116]*kernel[1]+tmp[5117]*kernel[2]+tmp[5215]*kernel[3]+tmp[5216]*kernel[4]+tmp[5217]*kernel[5]+tmp[5315]*kernel[6]+tmp[5316]*kernel[7]+tmp[5317]*kernel[8];
				ans[5217]<=tmp[5116]*kernel[0]+tmp[5117]*kernel[1]+tmp[5118]*kernel[2]+tmp[5216]*kernel[3]+tmp[5217]*kernel[4]+tmp[5218]*kernel[5]+tmp[5316]*kernel[6]+tmp[5317]*kernel[7]+tmp[5318]*kernel[8];
				ans[5218]<=tmp[5117]*kernel[0]+tmp[5118]*kernel[1]+tmp[5119]*kernel[2]+tmp[5217]*kernel[3]+tmp[5218]*kernel[4]+tmp[5219]*kernel[5]+tmp[5317]*kernel[6]+tmp[5318]*kernel[7]+tmp[5319]*kernel[8];
				ans[5219]<=tmp[5118]*kernel[0]+tmp[5119]*kernel[1]+tmp[5120]*kernel[2]+tmp[5218]*kernel[3]+tmp[5219]*kernel[4]+tmp[5220]*kernel[5]+tmp[5318]*kernel[6]+tmp[5319]*kernel[7]+tmp[5320]*kernel[8];
				ans[5220]<=tmp[5119]*kernel[0]+tmp[5120]*kernel[1]+tmp[5121]*kernel[2]+tmp[5219]*kernel[3]+tmp[5220]*kernel[4]+tmp[5221]*kernel[5]+tmp[5319]*kernel[6]+tmp[5320]*kernel[7]+tmp[5321]*kernel[8];
				ans[5221]<=tmp[5120]*kernel[0]+tmp[5121]*kernel[1]+tmp[5122]*kernel[2]+tmp[5220]*kernel[3]+tmp[5221]*kernel[4]+tmp[5222]*kernel[5]+tmp[5320]*kernel[6]+tmp[5321]*kernel[7]+tmp[5322]*kernel[8];
				ans[5222]<=tmp[5121]*kernel[0]+tmp[5122]*kernel[1]+tmp[5123]*kernel[2]+tmp[5221]*kernel[3]+tmp[5222]*kernel[4]+tmp[5223]*kernel[5]+tmp[5321]*kernel[6]+tmp[5322]*kernel[7]+tmp[5323]*kernel[8];
				ans[5223]<=tmp[5122]*kernel[0]+tmp[5123]*kernel[1]+tmp[5124]*kernel[2]+tmp[5222]*kernel[3]+tmp[5223]*kernel[4]+tmp[5224]*kernel[5]+tmp[5322]*kernel[6]+tmp[5323]*kernel[7]+tmp[5324]*kernel[8];
				ans[5224]<=tmp[5123]*kernel[0]+tmp[5124]*kernel[1]+tmp[5125]*kernel[2]+tmp[5223]*kernel[3]+tmp[5224]*kernel[4]+tmp[5225]*kernel[5]+tmp[5323]*kernel[6]+tmp[5324]*kernel[7]+tmp[5325]*kernel[8];
				ans[5225]<=tmp[5124]*kernel[0]+tmp[5125]*kernel[1]+tmp[5126]*kernel[2]+tmp[5224]*kernel[3]+tmp[5225]*kernel[4]+tmp[5226]*kernel[5]+tmp[5324]*kernel[6]+tmp[5325]*kernel[7]+tmp[5326]*kernel[8];
				ans[5226]<=tmp[5125]*kernel[0]+tmp[5126]*kernel[1]+tmp[5127]*kernel[2]+tmp[5225]*kernel[3]+tmp[5226]*kernel[4]+tmp[5227]*kernel[5]+tmp[5325]*kernel[6]+tmp[5326]*kernel[7]+tmp[5327]*kernel[8];
				ans[5227]<=tmp[5126]*kernel[0]+tmp[5127]*kernel[1]+tmp[5128]*kernel[2]+tmp[5226]*kernel[3]+tmp[5227]*kernel[4]+tmp[5228]*kernel[5]+tmp[5326]*kernel[6]+tmp[5327]*kernel[7]+tmp[5328]*kernel[8];
				ans[5228]<=tmp[5127]*kernel[0]+tmp[5128]*kernel[1]+tmp[5129]*kernel[2]+tmp[5227]*kernel[3]+tmp[5228]*kernel[4]+tmp[5229]*kernel[5]+tmp[5327]*kernel[6]+tmp[5328]*kernel[7]+tmp[5329]*kernel[8];
				ans[5229]<=tmp[5128]*kernel[0]+tmp[5129]*kernel[1]+tmp[5130]*kernel[2]+tmp[5228]*kernel[3]+tmp[5229]*kernel[4]+tmp[5230]*kernel[5]+tmp[5328]*kernel[6]+tmp[5329]*kernel[7]+tmp[5330]*kernel[8];
				ans[5230]<=tmp[5129]*kernel[0]+tmp[5130]*kernel[1]+tmp[5131]*kernel[2]+tmp[5229]*kernel[3]+tmp[5230]*kernel[4]+tmp[5231]*kernel[5]+tmp[5329]*kernel[6]+tmp[5330]*kernel[7]+tmp[5331]*kernel[8];
				ans[5231]<=tmp[5130]*kernel[0]+tmp[5131]*kernel[1]+tmp[5132]*kernel[2]+tmp[5230]*kernel[3]+tmp[5231]*kernel[4]+tmp[5232]*kernel[5]+tmp[5330]*kernel[6]+tmp[5331]*kernel[7]+tmp[5332]*kernel[8];
				ans[5232]<=tmp[5131]*kernel[0]+tmp[5132]*kernel[1]+tmp[5133]*kernel[2]+tmp[5231]*kernel[3]+tmp[5232]*kernel[4]+tmp[5233]*kernel[5]+tmp[5331]*kernel[6]+tmp[5332]*kernel[7]+tmp[5333]*kernel[8];
				ans[5233]<=tmp[5132]*kernel[0]+tmp[5133]*kernel[1]+tmp[5134]*kernel[2]+tmp[5232]*kernel[3]+tmp[5233]*kernel[4]+tmp[5234]*kernel[5]+tmp[5332]*kernel[6]+tmp[5333]*kernel[7]+tmp[5334]*kernel[8];
				ans[5234]<=tmp[5133]*kernel[0]+tmp[5134]*kernel[1]+tmp[5135]*kernel[2]+tmp[5233]*kernel[3]+tmp[5234]*kernel[4]+tmp[5235]*kernel[5]+tmp[5333]*kernel[6]+tmp[5334]*kernel[7]+tmp[5335]*kernel[8];
				ans[5235]<=tmp[5134]*kernel[0]+tmp[5135]*kernel[1]+tmp[5136]*kernel[2]+tmp[5234]*kernel[3]+tmp[5235]*kernel[4]+tmp[5236]*kernel[5]+tmp[5334]*kernel[6]+tmp[5335]*kernel[7]+tmp[5336]*kernel[8];
				ans[5236]<=tmp[5135]*kernel[0]+tmp[5136]*kernel[1]+tmp[5137]*kernel[2]+tmp[5235]*kernel[3]+tmp[5236]*kernel[4]+tmp[5237]*kernel[5]+tmp[5335]*kernel[6]+tmp[5336]*kernel[7]+tmp[5337]*kernel[8];
				ans[5237]<=tmp[5136]*kernel[0]+tmp[5137]*kernel[1]+tmp[5138]*kernel[2]+tmp[5236]*kernel[3]+tmp[5237]*kernel[4]+tmp[5238]*kernel[5]+tmp[5336]*kernel[6]+tmp[5337]*kernel[7]+tmp[5338]*kernel[8];
				ans[5238]<=tmp[5137]*kernel[0]+tmp[5138]*kernel[1]+tmp[5139]*kernel[2]+tmp[5237]*kernel[3]+tmp[5238]*kernel[4]+tmp[5239]*kernel[5]+tmp[5337]*kernel[6]+tmp[5338]*kernel[7]+tmp[5339]*kernel[8];
				ans[5239]<=tmp[5138]*kernel[0]+tmp[5139]*kernel[1]+tmp[5140]*kernel[2]+tmp[5238]*kernel[3]+tmp[5239]*kernel[4]+tmp[5240]*kernel[5]+tmp[5338]*kernel[6]+tmp[5339]*kernel[7]+tmp[5340]*kernel[8];
				ans[5240]<=tmp[5139]*kernel[0]+tmp[5140]*kernel[1]+tmp[5141]*kernel[2]+tmp[5239]*kernel[3]+tmp[5240]*kernel[4]+tmp[5241]*kernel[5]+tmp[5339]*kernel[6]+tmp[5340]*kernel[7]+tmp[5341]*kernel[8];
				ans[5241]<=tmp[5140]*kernel[0]+tmp[5141]*kernel[1]+tmp[5142]*kernel[2]+tmp[5240]*kernel[3]+tmp[5241]*kernel[4]+tmp[5242]*kernel[5]+tmp[5340]*kernel[6]+tmp[5341]*kernel[7]+tmp[5342]*kernel[8];
				ans[5242]<=tmp[5141]*kernel[0]+tmp[5142]*kernel[1]+tmp[5143]*kernel[2]+tmp[5241]*kernel[3]+tmp[5242]*kernel[4]+tmp[5243]*kernel[5]+tmp[5341]*kernel[6]+tmp[5342]*kernel[7]+tmp[5343]*kernel[8];
				ans[5243]<=tmp[5142]*kernel[0]+tmp[5143]*kernel[1]+tmp[5144]*kernel[2]+tmp[5242]*kernel[3]+tmp[5243]*kernel[4]+tmp[5244]*kernel[5]+tmp[5342]*kernel[6]+tmp[5343]*kernel[7]+tmp[5344]*kernel[8];
				ans[5244]<=tmp[5143]*kernel[0]+tmp[5144]*kernel[1]+tmp[5145]*kernel[2]+tmp[5243]*kernel[3]+tmp[5244]*kernel[4]+tmp[5245]*kernel[5]+tmp[5343]*kernel[6]+tmp[5344]*kernel[7]+tmp[5345]*kernel[8];
				ans[5245]<=tmp[5144]*kernel[0]+tmp[5145]*kernel[1]+tmp[5146]*kernel[2]+tmp[5244]*kernel[3]+tmp[5245]*kernel[4]+tmp[5246]*kernel[5]+tmp[5344]*kernel[6]+tmp[5345]*kernel[7]+tmp[5346]*kernel[8];
				ans[5246]<=tmp[5145]*kernel[0]+tmp[5146]*kernel[1]+tmp[5147]*kernel[2]+tmp[5245]*kernel[3]+tmp[5246]*kernel[4]+tmp[5247]*kernel[5]+tmp[5345]*kernel[6]+tmp[5346]*kernel[7]+tmp[5347]*kernel[8];
				ans[5247]<=tmp[5146]*kernel[0]+tmp[5147]*kernel[1]+tmp[5148]*kernel[2]+tmp[5246]*kernel[3]+tmp[5247]*kernel[4]+tmp[5248]*kernel[5]+tmp[5346]*kernel[6]+tmp[5347]*kernel[7]+tmp[5348]*kernel[8];
				ans[5248]<=tmp[5147]*kernel[0]+tmp[5148]*kernel[1]+tmp[5149]*kernel[2]+tmp[5247]*kernel[3]+tmp[5248]*kernel[4]+tmp[5249]*kernel[5]+tmp[5347]*kernel[6]+tmp[5348]*kernel[7]+tmp[5349]*kernel[8];
				ans[5249]<=tmp[5148]*kernel[0]+tmp[5149]*kernel[1]+tmp[5150]*kernel[2]+tmp[5248]*kernel[3]+tmp[5249]*kernel[4]+tmp[5250]*kernel[5]+tmp[5348]*kernel[6]+tmp[5349]*kernel[7]+tmp[5350]*kernel[8];
				ans[5250]<=tmp[5149]*kernel[0]+tmp[5150]*kernel[1]+tmp[5151]*kernel[2]+tmp[5249]*kernel[3]+tmp[5250]*kernel[4]+tmp[5251]*kernel[5]+tmp[5349]*kernel[6]+tmp[5350]*kernel[7]+tmp[5351]*kernel[8];
				ans[5251]<=tmp[5150]*kernel[0]+tmp[5151]*kernel[1]+tmp[5152]*kernel[2]+tmp[5250]*kernel[3]+tmp[5251]*kernel[4]+tmp[5252]*kernel[5]+tmp[5350]*kernel[6]+tmp[5351]*kernel[7]+tmp[5352]*kernel[8];
				ans[5252]<=tmp[5151]*kernel[0]+tmp[5152]*kernel[1]+tmp[5153]*kernel[2]+tmp[5251]*kernel[3]+tmp[5252]*kernel[4]+tmp[5253]*kernel[5]+tmp[5351]*kernel[6]+tmp[5352]*kernel[7]+tmp[5353]*kernel[8];
				ans[5253]<=tmp[5152]*kernel[0]+tmp[5153]*kernel[1]+tmp[5154]*kernel[2]+tmp[5252]*kernel[3]+tmp[5253]*kernel[4]+tmp[5254]*kernel[5]+tmp[5352]*kernel[6]+tmp[5353]*kernel[7]+tmp[5354]*kernel[8];
				ans[5254]<=tmp[5153]*kernel[0]+tmp[5154]*kernel[1]+tmp[5155]*kernel[2]+tmp[5253]*kernel[3]+tmp[5254]*kernel[4]+tmp[5255]*kernel[5]+tmp[5353]*kernel[6]+tmp[5354]*kernel[7]+tmp[5355]*kernel[8];
				ans[5255]<=tmp[5154]*kernel[0]+tmp[5155]*kernel[1]+tmp[5156]*kernel[2]+tmp[5254]*kernel[3]+tmp[5255]*kernel[4]+tmp[5256]*kernel[5]+tmp[5354]*kernel[6]+tmp[5355]*kernel[7]+tmp[5356]*kernel[8];
				ans[5256]<=tmp[5155]*kernel[0]+tmp[5156]*kernel[1]+tmp[5157]*kernel[2]+tmp[5255]*kernel[3]+tmp[5256]*kernel[4]+tmp[5257]*kernel[5]+tmp[5355]*kernel[6]+tmp[5356]*kernel[7]+tmp[5357]*kernel[8];
				ans[5257]<=tmp[5156]*kernel[0]+tmp[5157]*kernel[1]+tmp[5158]*kernel[2]+tmp[5256]*kernel[3]+tmp[5257]*kernel[4]+tmp[5258]*kernel[5]+tmp[5356]*kernel[6]+tmp[5357]*kernel[7]+tmp[5358]*kernel[8];
				ans[5258]<=tmp[5157]*kernel[0]+tmp[5158]*kernel[1]+tmp[5159]*kernel[2]+tmp[5257]*kernel[3]+tmp[5258]*kernel[4]+tmp[5259]*kernel[5]+tmp[5357]*kernel[6]+tmp[5358]*kernel[7]+tmp[5359]*kernel[8];
				ans[5259]<=tmp[5158]*kernel[0]+tmp[5159]*kernel[1]+tmp[5160]*kernel[2]+tmp[5258]*kernel[3]+tmp[5259]*kernel[4]+tmp[5260]*kernel[5]+tmp[5358]*kernel[6]+tmp[5359]*kernel[7]+tmp[5360]*kernel[8];
				ans[5260]<=tmp[5159]*kernel[0]+tmp[5160]*kernel[1]+tmp[5161]*kernel[2]+tmp[5259]*kernel[3]+tmp[5260]*kernel[4]+tmp[5261]*kernel[5]+tmp[5359]*kernel[6]+tmp[5360]*kernel[7]+tmp[5361]*kernel[8];
				ans[5261]<=tmp[5160]*kernel[0]+tmp[5161]*kernel[1]+tmp[5162]*kernel[2]+tmp[5260]*kernel[3]+tmp[5261]*kernel[4]+tmp[5262]*kernel[5]+tmp[5360]*kernel[6]+tmp[5361]*kernel[7]+tmp[5362]*kernel[8];
				ans[5262]<=tmp[5161]*kernel[0]+tmp[5162]*kernel[1]+tmp[5163]*kernel[2]+tmp[5261]*kernel[3]+tmp[5262]*kernel[4]+tmp[5263]*kernel[5]+tmp[5361]*kernel[6]+tmp[5362]*kernel[7]+tmp[5363]*kernel[8];
				ans[5263]<=tmp[5162]*kernel[0]+tmp[5163]*kernel[1]+tmp[5164]*kernel[2]+tmp[5262]*kernel[3]+tmp[5263]*kernel[4]+tmp[5264]*kernel[5]+tmp[5362]*kernel[6]+tmp[5363]*kernel[7]+tmp[5364]*kernel[8];
				ans[5264]<=tmp[5163]*kernel[0]+tmp[5164]*kernel[1]+tmp[5165]*kernel[2]+tmp[5263]*kernel[3]+tmp[5264]*kernel[4]+tmp[5265]*kernel[5]+tmp[5363]*kernel[6]+tmp[5364]*kernel[7]+tmp[5365]*kernel[8];
				ans[5265]<=tmp[5164]*kernel[0]+tmp[5165]*kernel[1]+tmp[5166]*kernel[2]+tmp[5264]*kernel[3]+tmp[5265]*kernel[4]+tmp[5266]*kernel[5]+tmp[5364]*kernel[6]+tmp[5365]*kernel[7]+tmp[5366]*kernel[8];
				ans[5266]<=tmp[5165]*kernel[0]+tmp[5166]*kernel[1]+tmp[5167]*kernel[2]+tmp[5265]*kernel[3]+tmp[5266]*kernel[4]+tmp[5267]*kernel[5]+tmp[5365]*kernel[6]+tmp[5366]*kernel[7]+tmp[5367]*kernel[8];
				ans[5267]<=tmp[5166]*kernel[0]+tmp[5167]*kernel[1]+tmp[5168]*kernel[2]+tmp[5266]*kernel[3]+tmp[5267]*kernel[4]+tmp[5268]*kernel[5]+tmp[5366]*kernel[6]+tmp[5367]*kernel[7]+tmp[5368]*kernel[8];
				ans[5268]<=tmp[5167]*kernel[0]+tmp[5168]*kernel[1]+tmp[5169]*kernel[2]+tmp[5267]*kernel[3]+tmp[5268]*kernel[4]+tmp[5269]*kernel[5]+tmp[5367]*kernel[6]+tmp[5368]*kernel[7]+tmp[5369]*kernel[8];
				ans[5269]<=tmp[5168]*kernel[0]+tmp[5169]*kernel[1]+tmp[5170]*kernel[2]+tmp[5268]*kernel[3]+tmp[5269]*kernel[4]+tmp[5270]*kernel[5]+tmp[5368]*kernel[6]+tmp[5369]*kernel[7]+tmp[5370]*kernel[8];
				ans[5270]<=tmp[5169]*kernel[0]+tmp[5170]*kernel[1]+tmp[5171]*kernel[2]+tmp[5269]*kernel[3]+tmp[5270]*kernel[4]+tmp[5271]*kernel[5]+tmp[5369]*kernel[6]+tmp[5370]*kernel[7]+tmp[5371]*kernel[8];
				ans[5271]<=tmp[5170]*kernel[0]+tmp[5171]*kernel[1]+tmp[5172]*kernel[2]+tmp[5270]*kernel[3]+tmp[5271]*kernel[4]+tmp[5272]*kernel[5]+tmp[5370]*kernel[6]+tmp[5371]*kernel[7]+tmp[5372]*kernel[8];
				ans[5272]<=tmp[5171]*kernel[0]+tmp[5172]*kernel[1]+tmp[5173]*kernel[2]+tmp[5271]*kernel[3]+tmp[5272]*kernel[4]+tmp[5273]*kernel[5]+tmp[5371]*kernel[6]+tmp[5372]*kernel[7]+tmp[5373]*kernel[8];
				ans[5273]<=tmp[5172]*kernel[0]+tmp[5173]*kernel[1]+tmp[5174]*kernel[2]+tmp[5272]*kernel[3]+tmp[5273]*kernel[4]+tmp[5274]*kernel[5]+tmp[5372]*kernel[6]+tmp[5373]*kernel[7]+tmp[5374]*kernel[8];
				ans[5274]<=tmp[5173]*kernel[0]+tmp[5174]*kernel[1]+tmp[5175]*kernel[2]+tmp[5273]*kernel[3]+tmp[5274]*kernel[4]+tmp[5275]*kernel[5]+tmp[5373]*kernel[6]+tmp[5374]*kernel[7]+tmp[5375]*kernel[8];
				ans[5275]<=tmp[5174]*kernel[0]+tmp[5175]*kernel[1]+tmp[5176]*kernel[2]+tmp[5274]*kernel[3]+tmp[5275]*kernel[4]+tmp[5276]*kernel[5]+tmp[5374]*kernel[6]+tmp[5375]*kernel[7]+tmp[5376]*kernel[8];
				ans[5276]<=tmp[5175]*kernel[0]+tmp[5176]*kernel[1]+tmp[5177]*kernel[2]+tmp[5275]*kernel[3]+tmp[5276]*kernel[4]+tmp[5277]*kernel[5]+tmp[5375]*kernel[6]+tmp[5376]*kernel[7]+tmp[5377]*kernel[8];
				ans[5277]<=tmp[5176]*kernel[0]+tmp[5177]*kernel[1]+tmp[5178]*kernel[2]+tmp[5276]*kernel[3]+tmp[5277]*kernel[4]+tmp[5278]*kernel[5]+tmp[5376]*kernel[6]+tmp[5377]*kernel[7]+tmp[5378]*kernel[8];
				ans[5278]<=tmp[5177]*kernel[0]+tmp[5178]*kernel[1]+tmp[5179]*kernel[2]+tmp[5277]*kernel[3]+tmp[5278]*kernel[4]+tmp[5279]*kernel[5]+tmp[5377]*kernel[6]+tmp[5378]*kernel[7]+tmp[5379]*kernel[8];
				ans[5279]<=tmp[5178]*kernel[0]+tmp[5179]*kernel[1]+tmp[5180]*kernel[2]+tmp[5278]*kernel[3]+tmp[5279]*kernel[4]+tmp[5280]*kernel[5]+tmp[5378]*kernel[6]+tmp[5379]*kernel[7]+tmp[5380]*kernel[8];
				ans[5280]<=tmp[5179]*kernel[0]+tmp[5180]*kernel[1]+tmp[5181]*kernel[2]+tmp[5279]*kernel[3]+tmp[5280]*kernel[4]+tmp[5281]*kernel[5]+tmp[5379]*kernel[6]+tmp[5380]*kernel[7]+tmp[5381]*kernel[8];
				ans[5281]<=tmp[5180]*kernel[0]+tmp[5181]*kernel[1]+tmp[5182]*kernel[2]+tmp[5280]*kernel[3]+tmp[5281]*kernel[4]+tmp[5282]*kernel[5]+tmp[5380]*kernel[6]+tmp[5381]*kernel[7]+tmp[5382]*kernel[8];
				ans[5282]<=tmp[5181]*kernel[0]+tmp[5182]*kernel[1]+tmp[5183]*kernel[2]+tmp[5281]*kernel[3]+tmp[5282]*kernel[4]+tmp[5283]*kernel[5]+tmp[5381]*kernel[6]+tmp[5382]*kernel[7]+tmp[5383]*kernel[8];
				ans[5283]<=tmp[5182]*kernel[0]+tmp[5183]*kernel[1]+tmp[5184]*kernel[2]+tmp[5282]*kernel[3]+tmp[5283]*kernel[4]+tmp[5284]*kernel[5]+tmp[5382]*kernel[6]+tmp[5383]*kernel[7]+tmp[5384]*kernel[8];
				ans[5284]<=tmp[5183]*kernel[0]+tmp[5184]*kernel[1]+tmp[5185]*kernel[2]+tmp[5283]*kernel[3]+tmp[5284]*kernel[4]+tmp[5285]*kernel[5]+tmp[5383]*kernel[6]+tmp[5384]*kernel[7]+tmp[5385]*kernel[8];
				ans[5285]<=tmp[5184]*kernel[0]+tmp[5185]*kernel[1]+tmp[5186]*kernel[2]+tmp[5284]*kernel[3]+tmp[5285]*kernel[4]+tmp[5286]*kernel[5]+tmp[5384]*kernel[6]+tmp[5385]*kernel[7]+tmp[5386]*kernel[8];
				ans[5286]<=tmp[5185]*kernel[0]+tmp[5186]*kernel[1]+tmp[5187]*kernel[2]+tmp[5285]*kernel[3]+tmp[5286]*kernel[4]+tmp[5287]*kernel[5]+tmp[5385]*kernel[6]+tmp[5386]*kernel[7]+tmp[5387]*kernel[8];
				ans[5287]<=tmp[5186]*kernel[0]+tmp[5187]*kernel[1]+tmp[5188]*kernel[2]+tmp[5286]*kernel[3]+tmp[5287]*kernel[4]+tmp[5288]*kernel[5]+tmp[5386]*kernel[6]+tmp[5387]*kernel[7]+tmp[5388]*kernel[8];
				ans[5288]<=tmp[5187]*kernel[0]+tmp[5188]*kernel[1]+tmp[5189]*kernel[2]+tmp[5287]*kernel[3]+tmp[5288]*kernel[4]+tmp[5289]*kernel[5]+tmp[5387]*kernel[6]+tmp[5388]*kernel[7]+tmp[5389]*kernel[8];
				ans[5289]<=tmp[5188]*kernel[0]+tmp[5189]*kernel[1]+tmp[5190]*kernel[2]+tmp[5288]*kernel[3]+tmp[5289]*kernel[4]+tmp[5290]*kernel[5]+tmp[5388]*kernel[6]+tmp[5389]*kernel[7]+tmp[5390]*kernel[8];
				ans[5290]<=tmp[5189]*kernel[0]+tmp[5190]*kernel[1]+tmp[5191]*kernel[2]+tmp[5289]*kernel[3]+tmp[5290]*kernel[4]+tmp[5291]*kernel[5]+tmp[5389]*kernel[6]+tmp[5390]*kernel[7]+tmp[5391]*kernel[8];
				ans[5291]<=tmp[5190]*kernel[0]+tmp[5191]*kernel[1]+tmp[5192]*kernel[2]+tmp[5290]*kernel[3]+tmp[5291]*kernel[4]+tmp[5292]*kernel[5]+tmp[5390]*kernel[6]+tmp[5391]*kernel[7]+tmp[5392]*kernel[8];
				ans[5292]<=tmp[5191]*kernel[0]+tmp[5192]*kernel[1]+tmp[5193]*kernel[2]+tmp[5291]*kernel[3]+tmp[5292]*kernel[4]+tmp[5293]*kernel[5]+tmp[5391]*kernel[6]+tmp[5392]*kernel[7]+tmp[5393]*kernel[8];
				ans[5293]<=tmp[5192]*kernel[0]+tmp[5193]*kernel[1]+tmp[5194]*kernel[2]+tmp[5292]*kernel[3]+tmp[5293]*kernel[4]+tmp[5294]*kernel[5]+tmp[5392]*kernel[6]+tmp[5393]*kernel[7]+tmp[5394]*kernel[8];
				ans[5294]<=tmp[5193]*kernel[0]+tmp[5194]*kernel[1]+tmp[5195]*kernel[2]+tmp[5293]*kernel[3]+tmp[5294]*kernel[4]+tmp[5295]*kernel[5]+tmp[5393]*kernel[6]+tmp[5394]*kernel[7]+tmp[5395]*kernel[8];
				ans[5295]<=tmp[5194]*kernel[0]+tmp[5195]*kernel[1]+tmp[5196]*kernel[2]+tmp[5294]*kernel[3]+tmp[5295]*kernel[4]+tmp[5296]*kernel[5]+tmp[5394]*kernel[6]+tmp[5395]*kernel[7]+tmp[5396]*kernel[8];
				ans[5296]<=tmp[5195]*kernel[0]+tmp[5196]*kernel[1]+tmp[5197]*kernel[2]+tmp[5295]*kernel[3]+tmp[5296]*kernel[4]+tmp[5297]*kernel[5]+tmp[5395]*kernel[6]+tmp[5396]*kernel[7]+tmp[5397]*kernel[8];
				ans[5297]<=tmp[5196]*kernel[0]+tmp[5197]*kernel[1]+tmp[5198]*kernel[2]+tmp[5296]*kernel[3]+tmp[5297]*kernel[4]+tmp[5298]*kernel[5]+tmp[5396]*kernel[6]+tmp[5397]*kernel[7]+tmp[5398]*kernel[8];
				ans[5298]<=tmp[5197]*kernel[0]+tmp[5198]*kernel[1]+tmp[5199]*kernel[2]+tmp[5297]*kernel[3]+tmp[5298]*kernel[4]+tmp[5299]*kernel[5]+tmp[5397]*kernel[6]+tmp[5398]*kernel[7]+tmp[5399]*kernel[8];
				ans[5299]<=tmp[5198]*kernel[0]+tmp[5199]*kernel[1]+tmp[5298]*kernel[3]+tmp[5299]*kernel[4]+tmp[5398]*kernel[6]+tmp[5399]*kernel[7];
				ans[5300]<=tmp[5200]*kernel[1]+tmp[5201]*kernel[2]+tmp[5300]*kernel[4]+tmp[5301]*kernel[5]+tmp[5400]*kernel[7]+tmp[5401]*kernel[8];
				ans[5301]<=tmp[5200]*kernel[0]+tmp[5201]*kernel[1]+tmp[5202]*kernel[2]+tmp[5300]*kernel[3]+tmp[5301]*kernel[4]+tmp[5302]*kernel[5]+tmp[5400]*kernel[6]+tmp[5401]*kernel[7]+tmp[5402]*kernel[8];
				ans[5302]<=tmp[5201]*kernel[0]+tmp[5202]*kernel[1]+tmp[5203]*kernel[2]+tmp[5301]*kernel[3]+tmp[5302]*kernel[4]+tmp[5303]*kernel[5]+tmp[5401]*kernel[6]+tmp[5402]*kernel[7]+tmp[5403]*kernel[8];
				ans[5303]<=tmp[5202]*kernel[0]+tmp[5203]*kernel[1]+tmp[5204]*kernel[2]+tmp[5302]*kernel[3]+tmp[5303]*kernel[4]+tmp[5304]*kernel[5]+tmp[5402]*kernel[6]+tmp[5403]*kernel[7]+tmp[5404]*kernel[8];
				ans[5304]<=tmp[5203]*kernel[0]+tmp[5204]*kernel[1]+tmp[5205]*kernel[2]+tmp[5303]*kernel[3]+tmp[5304]*kernel[4]+tmp[5305]*kernel[5]+tmp[5403]*kernel[6]+tmp[5404]*kernel[7]+tmp[5405]*kernel[8];
				ans[5305]<=tmp[5204]*kernel[0]+tmp[5205]*kernel[1]+tmp[5206]*kernel[2]+tmp[5304]*kernel[3]+tmp[5305]*kernel[4]+tmp[5306]*kernel[5]+tmp[5404]*kernel[6]+tmp[5405]*kernel[7]+tmp[5406]*kernel[8];
				ans[5306]<=tmp[5205]*kernel[0]+tmp[5206]*kernel[1]+tmp[5207]*kernel[2]+tmp[5305]*kernel[3]+tmp[5306]*kernel[4]+tmp[5307]*kernel[5]+tmp[5405]*kernel[6]+tmp[5406]*kernel[7]+tmp[5407]*kernel[8];
				ans[5307]<=tmp[5206]*kernel[0]+tmp[5207]*kernel[1]+tmp[5208]*kernel[2]+tmp[5306]*kernel[3]+tmp[5307]*kernel[4]+tmp[5308]*kernel[5]+tmp[5406]*kernel[6]+tmp[5407]*kernel[7]+tmp[5408]*kernel[8];
				ans[5308]<=tmp[5207]*kernel[0]+tmp[5208]*kernel[1]+tmp[5209]*kernel[2]+tmp[5307]*kernel[3]+tmp[5308]*kernel[4]+tmp[5309]*kernel[5]+tmp[5407]*kernel[6]+tmp[5408]*kernel[7]+tmp[5409]*kernel[8];
				ans[5309]<=tmp[5208]*kernel[0]+tmp[5209]*kernel[1]+tmp[5210]*kernel[2]+tmp[5308]*kernel[3]+tmp[5309]*kernel[4]+tmp[5310]*kernel[5]+tmp[5408]*kernel[6]+tmp[5409]*kernel[7]+tmp[5410]*kernel[8];
				ans[5310]<=tmp[5209]*kernel[0]+tmp[5210]*kernel[1]+tmp[5211]*kernel[2]+tmp[5309]*kernel[3]+tmp[5310]*kernel[4]+tmp[5311]*kernel[5]+tmp[5409]*kernel[6]+tmp[5410]*kernel[7]+tmp[5411]*kernel[8];
				ans[5311]<=tmp[5210]*kernel[0]+tmp[5211]*kernel[1]+tmp[5212]*kernel[2]+tmp[5310]*kernel[3]+tmp[5311]*kernel[4]+tmp[5312]*kernel[5]+tmp[5410]*kernel[6]+tmp[5411]*kernel[7]+tmp[5412]*kernel[8];
				ans[5312]<=tmp[5211]*kernel[0]+tmp[5212]*kernel[1]+tmp[5213]*kernel[2]+tmp[5311]*kernel[3]+tmp[5312]*kernel[4]+tmp[5313]*kernel[5]+tmp[5411]*kernel[6]+tmp[5412]*kernel[7]+tmp[5413]*kernel[8];
				ans[5313]<=tmp[5212]*kernel[0]+tmp[5213]*kernel[1]+tmp[5214]*kernel[2]+tmp[5312]*kernel[3]+tmp[5313]*kernel[4]+tmp[5314]*kernel[5]+tmp[5412]*kernel[6]+tmp[5413]*kernel[7]+tmp[5414]*kernel[8];
				ans[5314]<=tmp[5213]*kernel[0]+tmp[5214]*kernel[1]+tmp[5215]*kernel[2]+tmp[5313]*kernel[3]+tmp[5314]*kernel[4]+tmp[5315]*kernel[5]+tmp[5413]*kernel[6]+tmp[5414]*kernel[7]+tmp[5415]*kernel[8];
				ans[5315]<=tmp[5214]*kernel[0]+tmp[5215]*kernel[1]+tmp[5216]*kernel[2]+tmp[5314]*kernel[3]+tmp[5315]*kernel[4]+tmp[5316]*kernel[5]+tmp[5414]*kernel[6]+tmp[5415]*kernel[7]+tmp[5416]*kernel[8];
				ans[5316]<=tmp[5215]*kernel[0]+tmp[5216]*kernel[1]+tmp[5217]*kernel[2]+tmp[5315]*kernel[3]+tmp[5316]*kernel[4]+tmp[5317]*kernel[5]+tmp[5415]*kernel[6]+tmp[5416]*kernel[7]+tmp[5417]*kernel[8];
				ans[5317]<=tmp[5216]*kernel[0]+tmp[5217]*kernel[1]+tmp[5218]*kernel[2]+tmp[5316]*kernel[3]+tmp[5317]*kernel[4]+tmp[5318]*kernel[5]+tmp[5416]*kernel[6]+tmp[5417]*kernel[7]+tmp[5418]*kernel[8];
				ans[5318]<=tmp[5217]*kernel[0]+tmp[5218]*kernel[1]+tmp[5219]*kernel[2]+tmp[5317]*kernel[3]+tmp[5318]*kernel[4]+tmp[5319]*kernel[5]+tmp[5417]*kernel[6]+tmp[5418]*kernel[7]+tmp[5419]*kernel[8];
				ans[5319]<=tmp[5218]*kernel[0]+tmp[5219]*kernel[1]+tmp[5220]*kernel[2]+tmp[5318]*kernel[3]+tmp[5319]*kernel[4]+tmp[5320]*kernel[5]+tmp[5418]*kernel[6]+tmp[5419]*kernel[7]+tmp[5420]*kernel[8];
				ans[5320]<=tmp[5219]*kernel[0]+tmp[5220]*kernel[1]+tmp[5221]*kernel[2]+tmp[5319]*kernel[3]+tmp[5320]*kernel[4]+tmp[5321]*kernel[5]+tmp[5419]*kernel[6]+tmp[5420]*kernel[7]+tmp[5421]*kernel[8];
				ans[5321]<=tmp[5220]*kernel[0]+tmp[5221]*kernel[1]+tmp[5222]*kernel[2]+tmp[5320]*kernel[3]+tmp[5321]*kernel[4]+tmp[5322]*kernel[5]+tmp[5420]*kernel[6]+tmp[5421]*kernel[7]+tmp[5422]*kernel[8];
				ans[5322]<=tmp[5221]*kernel[0]+tmp[5222]*kernel[1]+tmp[5223]*kernel[2]+tmp[5321]*kernel[3]+tmp[5322]*kernel[4]+tmp[5323]*kernel[5]+tmp[5421]*kernel[6]+tmp[5422]*kernel[7]+tmp[5423]*kernel[8];
				ans[5323]<=tmp[5222]*kernel[0]+tmp[5223]*kernel[1]+tmp[5224]*kernel[2]+tmp[5322]*kernel[3]+tmp[5323]*kernel[4]+tmp[5324]*kernel[5]+tmp[5422]*kernel[6]+tmp[5423]*kernel[7]+tmp[5424]*kernel[8];
				ans[5324]<=tmp[5223]*kernel[0]+tmp[5224]*kernel[1]+tmp[5225]*kernel[2]+tmp[5323]*kernel[3]+tmp[5324]*kernel[4]+tmp[5325]*kernel[5]+tmp[5423]*kernel[6]+tmp[5424]*kernel[7]+tmp[5425]*kernel[8];
				ans[5325]<=tmp[5224]*kernel[0]+tmp[5225]*kernel[1]+tmp[5226]*kernel[2]+tmp[5324]*kernel[3]+tmp[5325]*kernel[4]+tmp[5326]*kernel[5]+tmp[5424]*kernel[6]+tmp[5425]*kernel[7]+tmp[5426]*kernel[8];
				ans[5326]<=tmp[5225]*kernel[0]+tmp[5226]*kernel[1]+tmp[5227]*kernel[2]+tmp[5325]*kernel[3]+tmp[5326]*kernel[4]+tmp[5327]*kernel[5]+tmp[5425]*kernel[6]+tmp[5426]*kernel[7]+tmp[5427]*kernel[8];
				ans[5327]<=tmp[5226]*kernel[0]+tmp[5227]*kernel[1]+tmp[5228]*kernel[2]+tmp[5326]*kernel[3]+tmp[5327]*kernel[4]+tmp[5328]*kernel[5]+tmp[5426]*kernel[6]+tmp[5427]*kernel[7]+tmp[5428]*kernel[8];
				ans[5328]<=tmp[5227]*kernel[0]+tmp[5228]*kernel[1]+tmp[5229]*kernel[2]+tmp[5327]*kernel[3]+tmp[5328]*kernel[4]+tmp[5329]*kernel[5]+tmp[5427]*kernel[6]+tmp[5428]*kernel[7]+tmp[5429]*kernel[8];
				ans[5329]<=tmp[5228]*kernel[0]+tmp[5229]*kernel[1]+tmp[5230]*kernel[2]+tmp[5328]*kernel[3]+tmp[5329]*kernel[4]+tmp[5330]*kernel[5]+tmp[5428]*kernel[6]+tmp[5429]*kernel[7]+tmp[5430]*kernel[8];
				ans[5330]<=tmp[5229]*kernel[0]+tmp[5230]*kernel[1]+tmp[5231]*kernel[2]+tmp[5329]*kernel[3]+tmp[5330]*kernel[4]+tmp[5331]*kernel[5]+tmp[5429]*kernel[6]+tmp[5430]*kernel[7]+tmp[5431]*kernel[8];
				ans[5331]<=tmp[5230]*kernel[0]+tmp[5231]*kernel[1]+tmp[5232]*kernel[2]+tmp[5330]*kernel[3]+tmp[5331]*kernel[4]+tmp[5332]*kernel[5]+tmp[5430]*kernel[6]+tmp[5431]*kernel[7]+tmp[5432]*kernel[8];
				ans[5332]<=tmp[5231]*kernel[0]+tmp[5232]*kernel[1]+tmp[5233]*kernel[2]+tmp[5331]*kernel[3]+tmp[5332]*kernel[4]+tmp[5333]*kernel[5]+tmp[5431]*kernel[6]+tmp[5432]*kernel[7]+tmp[5433]*kernel[8];
				ans[5333]<=tmp[5232]*kernel[0]+tmp[5233]*kernel[1]+tmp[5234]*kernel[2]+tmp[5332]*kernel[3]+tmp[5333]*kernel[4]+tmp[5334]*kernel[5]+tmp[5432]*kernel[6]+tmp[5433]*kernel[7]+tmp[5434]*kernel[8];
				ans[5334]<=tmp[5233]*kernel[0]+tmp[5234]*kernel[1]+tmp[5235]*kernel[2]+tmp[5333]*kernel[3]+tmp[5334]*kernel[4]+tmp[5335]*kernel[5]+tmp[5433]*kernel[6]+tmp[5434]*kernel[7]+tmp[5435]*kernel[8];
				ans[5335]<=tmp[5234]*kernel[0]+tmp[5235]*kernel[1]+tmp[5236]*kernel[2]+tmp[5334]*kernel[3]+tmp[5335]*kernel[4]+tmp[5336]*kernel[5]+tmp[5434]*kernel[6]+tmp[5435]*kernel[7]+tmp[5436]*kernel[8];
				ans[5336]<=tmp[5235]*kernel[0]+tmp[5236]*kernel[1]+tmp[5237]*kernel[2]+tmp[5335]*kernel[3]+tmp[5336]*kernel[4]+tmp[5337]*kernel[5]+tmp[5435]*kernel[6]+tmp[5436]*kernel[7]+tmp[5437]*kernel[8];
				ans[5337]<=tmp[5236]*kernel[0]+tmp[5237]*kernel[1]+tmp[5238]*kernel[2]+tmp[5336]*kernel[3]+tmp[5337]*kernel[4]+tmp[5338]*kernel[5]+tmp[5436]*kernel[6]+tmp[5437]*kernel[7]+tmp[5438]*kernel[8];
				ans[5338]<=tmp[5237]*kernel[0]+tmp[5238]*kernel[1]+tmp[5239]*kernel[2]+tmp[5337]*kernel[3]+tmp[5338]*kernel[4]+tmp[5339]*kernel[5]+tmp[5437]*kernel[6]+tmp[5438]*kernel[7]+tmp[5439]*kernel[8];
				ans[5339]<=tmp[5238]*kernel[0]+tmp[5239]*kernel[1]+tmp[5240]*kernel[2]+tmp[5338]*kernel[3]+tmp[5339]*kernel[4]+tmp[5340]*kernel[5]+tmp[5438]*kernel[6]+tmp[5439]*kernel[7]+tmp[5440]*kernel[8];
				ans[5340]<=tmp[5239]*kernel[0]+tmp[5240]*kernel[1]+tmp[5241]*kernel[2]+tmp[5339]*kernel[3]+tmp[5340]*kernel[4]+tmp[5341]*kernel[5]+tmp[5439]*kernel[6]+tmp[5440]*kernel[7]+tmp[5441]*kernel[8];
				ans[5341]<=tmp[5240]*kernel[0]+tmp[5241]*kernel[1]+tmp[5242]*kernel[2]+tmp[5340]*kernel[3]+tmp[5341]*kernel[4]+tmp[5342]*kernel[5]+tmp[5440]*kernel[6]+tmp[5441]*kernel[7]+tmp[5442]*kernel[8];
				ans[5342]<=tmp[5241]*kernel[0]+tmp[5242]*kernel[1]+tmp[5243]*kernel[2]+tmp[5341]*kernel[3]+tmp[5342]*kernel[4]+tmp[5343]*kernel[5]+tmp[5441]*kernel[6]+tmp[5442]*kernel[7]+tmp[5443]*kernel[8];
				ans[5343]<=tmp[5242]*kernel[0]+tmp[5243]*kernel[1]+tmp[5244]*kernel[2]+tmp[5342]*kernel[3]+tmp[5343]*kernel[4]+tmp[5344]*kernel[5]+tmp[5442]*kernel[6]+tmp[5443]*kernel[7]+tmp[5444]*kernel[8];
				ans[5344]<=tmp[5243]*kernel[0]+tmp[5244]*kernel[1]+tmp[5245]*kernel[2]+tmp[5343]*kernel[3]+tmp[5344]*kernel[4]+tmp[5345]*kernel[5]+tmp[5443]*kernel[6]+tmp[5444]*kernel[7]+tmp[5445]*kernel[8];
				ans[5345]<=tmp[5244]*kernel[0]+tmp[5245]*kernel[1]+tmp[5246]*kernel[2]+tmp[5344]*kernel[3]+tmp[5345]*kernel[4]+tmp[5346]*kernel[5]+tmp[5444]*kernel[6]+tmp[5445]*kernel[7]+tmp[5446]*kernel[8];
				ans[5346]<=tmp[5245]*kernel[0]+tmp[5246]*kernel[1]+tmp[5247]*kernel[2]+tmp[5345]*kernel[3]+tmp[5346]*kernel[4]+tmp[5347]*kernel[5]+tmp[5445]*kernel[6]+tmp[5446]*kernel[7]+tmp[5447]*kernel[8];
				ans[5347]<=tmp[5246]*kernel[0]+tmp[5247]*kernel[1]+tmp[5248]*kernel[2]+tmp[5346]*kernel[3]+tmp[5347]*kernel[4]+tmp[5348]*kernel[5]+tmp[5446]*kernel[6]+tmp[5447]*kernel[7]+tmp[5448]*kernel[8];
				ans[5348]<=tmp[5247]*kernel[0]+tmp[5248]*kernel[1]+tmp[5249]*kernel[2]+tmp[5347]*kernel[3]+tmp[5348]*kernel[4]+tmp[5349]*kernel[5]+tmp[5447]*kernel[6]+tmp[5448]*kernel[7]+tmp[5449]*kernel[8];
				ans[5349]<=tmp[5248]*kernel[0]+tmp[5249]*kernel[1]+tmp[5250]*kernel[2]+tmp[5348]*kernel[3]+tmp[5349]*kernel[4]+tmp[5350]*kernel[5]+tmp[5448]*kernel[6]+tmp[5449]*kernel[7]+tmp[5450]*kernel[8];
				ans[5350]<=tmp[5249]*kernel[0]+tmp[5250]*kernel[1]+tmp[5251]*kernel[2]+tmp[5349]*kernel[3]+tmp[5350]*kernel[4]+tmp[5351]*kernel[5]+tmp[5449]*kernel[6]+tmp[5450]*kernel[7]+tmp[5451]*kernel[8];
				ans[5351]<=tmp[5250]*kernel[0]+tmp[5251]*kernel[1]+tmp[5252]*kernel[2]+tmp[5350]*kernel[3]+tmp[5351]*kernel[4]+tmp[5352]*kernel[5]+tmp[5450]*kernel[6]+tmp[5451]*kernel[7]+tmp[5452]*kernel[8];
				ans[5352]<=tmp[5251]*kernel[0]+tmp[5252]*kernel[1]+tmp[5253]*kernel[2]+tmp[5351]*kernel[3]+tmp[5352]*kernel[4]+tmp[5353]*kernel[5]+tmp[5451]*kernel[6]+tmp[5452]*kernel[7]+tmp[5453]*kernel[8];
				ans[5353]<=tmp[5252]*kernel[0]+tmp[5253]*kernel[1]+tmp[5254]*kernel[2]+tmp[5352]*kernel[3]+tmp[5353]*kernel[4]+tmp[5354]*kernel[5]+tmp[5452]*kernel[6]+tmp[5453]*kernel[7]+tmp[5454]*kernel[8];
				ans[5354]<=tmp[5253]*kernel[0]+tmp[5254]*kernel[1]+tmp[5255]*kernel[2]+tmp[5353]*kernel[3]+tmp[5354]*kernel[4]+tmp[5355]*kernel[5]+tmp[5453]*kernel[6]+tmp[5454]*kernel[7]+tmp[5455]*kernel[8];
				ans[5355]<=tmp[5254]*kernel[0]+tmp[5255]*kernel[1]+tmp[5256]*kernel[2]+tmp[5354]*kernel[3]+tmp[5355]*kernel[4]+tmp[5356]*kernel[5]+tmp[5454]*kernel[6]+tmp[5455]*kernel[7]+tmp[5456]*kernel[8];
				ans[5356]<=tmp[5255]*kernel[0]+tmp[5256]*kernel[1]+tmp[5257]*kernel[2]+tmp[5355]*kernel[3]+tmp[5356]*kernel[4]+tmp[5357]*kernel[5]+tmp[5455]*kernel[6]+tmp[5456]*kernel[7]+tmp[5457]*kernel[8];
				ans[5357]<=tmp[5256]*kernel[0]+tmp[5257]*kernel[1]+tmp[5258]*kernel[2]+tmp[5356]*kernel[3]+tmp[5357]*kernel[4]+tmp[5358]*kernel[5]+tmp[5456]*kernel[6]+tmp[5457]*kernel[7]+tmp[5458]*kernel[8];
				ans[5358]<=tmp[5257]*kernel[0]+tmp[5258]*kernel[1]+tmp[5259]*kernel[2]+tmp[5357]*kernel[3]+tmp[5358]*kernel[4]+tmp[5359]*kernel[5]+tmp[5457]*kernel[6]+tmp[5458]*kernel[7]+tmp[5459]*kernel[8];
				ans[5359]<=tmp[5258]*kernel[0]+tmp[5259]*kernel[1]+tmp[5260]*kernel[2]+tmp[5358]*kernel[3]+tmp[5359]*kernel[4]+tmp[5360]*kernel[5]+tmp[5458]*kernel[6]+tmp[5459]*kernel[7]+tmp[5460]*kernel[8];
				ans[5360]<=tmp[5259]*kernel[0]+tmp[5260]*kernel[1]+tmp[5261]*kernel[2]+tmp[5359]*kernel[3]+tmp[5360]*kernel[4]+tmp[5361]*kernel[5]+tmp[5459]*kernel[6]+tmp[5460]*kernel[7]+tmp[5461]*kernel[8];
				ans[5361]<=tmp[5260]*kernel[0]+tmp[5261]*kernel[1]+tmp[5262]*kernel[2]+tmp[5360]*kernel[3]+tmp[5361]*kernel[4]+tmp[5362]*kernel[5]+tmp[5460]*kernel[6]+tmp[5461]*kernel[7]+tmp[5462]*kernel[8];
				ans[5362]<=tmp[5261]*kernel[0]+tmp[5262]*kernel[1]+tmp[5263]*kernel[2]+tmp[5361]*kernel[3]+tmp[5362]*kernel[4]+tmp[5363]*kernel[5]+tmp[5461]*kernel[6]+tmp[5462]*kernel[7]+tmp[5463]*kernel[8];
				ans[5363]<=tmp[5262]*kernel[0]+tmp[5263]*kernel[1]+tmp[5264]*kernel[2]+tmp[5362]*kernel[3]+tmp[5363]*kernel[4]+tmp[5364]*kernel[5]+tmp[5462]*kernel[6]+tmp[5463]*kernel[7]+tmp[5464]*kernel[8];
				ans[5364]<=tmp[5263]*kernel[0]+tmp[5264]*kernel[1]+tmp[5265]*kernel[2]+tmp[5363]*kernel[3]+tmp[5364]*kernel[4]+tmp[5365]*kernel[5]+tmp[5463]*kernel[6]+tmp[5464]*kernel[7]+tmp[5465]*kernel[8];
				ans[5365]<=tmp[5264]*kernel[0]+tmp[5265]*kernel[1]+tmp[5266]*kernel[2]+tmp[5364]*kernel[3]+tmp[5365]*kernel[4]+tmp[5366]*kernel[5]+tmp[5464]*kernel[6]+tmp[5465]*kernel[7]+tmp[5466]*kernel[8];
				ans[5366]<=tmp[5265]*kernel[0]+tmp[5266]*kernel[1]+tmp[5267]*kernel[2]+tmp[5365]*kernel[3]+tmp[5366]*kernel[4]+tmp[5367]*kernel[5]+tmp[5465]*kernel[6]+tmp[5466]*kernel[7]+tmp[5467]*kernel[8];
				ans[5367]<=tmp[5266]*kernel[0]+tmp[5267]*kernel[1]+tmp[5268]*kernel[2]+tmp[5366]*kernel[3]+tmp[5367]*kernel[4]+tmp[5368]*kernel[5]+tmp[5466]*kernel[6]+tmp[5467]*kernel[7]+tmp[5468]*kernel[8];
				ans[5368]<=tmp[5267]*kernel[0]+tmp[5268]*kernel[1]+tmp[5269]*kernel[2]+tmp[5367]*kernel[3]+tmp[5368]*kernel[4]+tmp[5369]*kernel[5]+tmp[5467]*kernel[6]+tmp[5468]*kernel[7]+tmp[5469]*kernel[8];
				ans[5369]<=tmp[5268]*kernel[0]+tmp[5269]*kernel[1]+tmp[5270]*kernel[2]+tmp[5368]*kernel[3]+tmp[5369]*kernel[4]+tmp[5370]*kernel[5]+tmp[5468]*kernel[6]+tmp[5469]*kernel[7]+tmp[5470]*kernel[8];
				ans[5370]<=tmp[5269]*kernel[0]+tmp[5270]*kernel[1]+tmp[5271]*kernel[2]+tmp[5369]*kernel[3]+tmp[5370]*kernel[4]+tmp[5371]*kernel[5]+tmp[5469]*kernel[6]+tmp[5470]*kernel[7]+tmp[5471]*kernel[8];
				ans[5371]<=tmp[5270]*kernel[0]+tmp[5271]*kernel[1]+tmp[5272]*kernel[2]+tmp[5370]*kernel[3]+tmp[5371]*kernel[4]+tmp[5372]*kernel[5]+tmp[5470]*kernel[6]+tmp[5471]*kernel[7]+tmp[5472]*kernel[8];
				ans[5372]<=tmp[5271]*kernel[0]+tmp[5272]*kernel[1]+tmp[5273]*kernel[2]+tmp[5371]*kernel[3]+tmp[5372]*kernel[4]+tmp[5373]*kernel[5]+tmp[5471]*kernel[6]+tmp[5472]*kernel[7]+tmp[5473]*kernel[8];
				ans[5373]<=tmp[5272]*kernel[0]+tmp[5273]*kernel[1]+tmp[5274]*kernel[2]+tmp[5372]*kernel[3]+tmp[5373]*kernel[4]+tmp[5374]*kernel[5]+tmp[5472]*kernel[6]+tmp[5473]*kernel[7]+tmp[5474]*kernel[8];
				ans[5374]<=tmp[5273]*kernel[0]+tmp[5274]*kernel[1]+tmp[5275]*kernel[2]+tmp[5373]*kernel[3]+tmp[5374]*kernel[4]+tmp[5375]*kernel[5]+tmp[5473]*kernel[6]+tmp[5474]*kernel[7]+tmp[5475]*kernel[8];
				ans[5375]<=tmp[5274]*kernel[0]+tmp[5275]*kernel[1]+tmp[5276]*kernel[2]+tmp[5374]*kernel[3]+tmp[5375]*kernel[4]+tmp[5376]*kernel[5]+tmp[5474]*kernel[6]+tmp[5475]*kernel[7]+tmp[5476]*kernel[8];
				ans[5376]<=tmp[5275]*kernel[0]+tmp[5276]*kernel[1]+tmp[5277]*kernel[2]+tmp[5375]*kernel[3]+tmp[5376]*kernel[4]+tmp[5377]*kernel[5]+tmp[5475]*kernel[6]+tmp[5476]*kernel[7]+tmp[5477]*kernel[8];
				ans[5377]<=tmp[5276]*kernel[0]+tmp[5277]*kernel[1]+tmp[5278]*kernel[2]+tmp[5376]*kernel[3]+tmp[5377]*kernel[4]+tmp[5378]*kernel[5]+tmp[5476]*kernel[6]+tmp[5477]*kernel[7]+tmp[5478]*kernel[8];
				ans[5378]<=tmp[5277]*kernel[0]+tmp[5278]*kernel[1]+tmp[5279]*kernel[2]+tmp[5377]*kernel[3]+tmp[5378]*kernel[4]+tmp[5379]*kernel[5]+tmp[5477]*kernel[6]+tmp[5478]*kernel[7]+tmp[5479]*kernel[8];
				ans[5379]<=tmp[5278]*kernel[0]+tmp[5279]*kernel[1]+tmp[5280]*kernel[2]+tmp[5378]*kernel[3]+tmp[5379]*kernel[4]+tmp[5380]*kernel[5]+tmp[5478]*kernel[6]+tmp[5479]*kernel[7]+tmp[5480]*kernel[8];
				ans[5380]<=tmp[5279]*kernel[0]+tmp[5280]*kernel[1]+tmp[5281]*kernel[2]+tmp[5379]*kernel[3]+tmp[5380]*kernel[4]+tmp[5381]*kernel[5]+tmp[5479]*kernel[6]+tmp[5480]*kernel[7]+tmp[5481]*kernel[8];
				ans[5381]<=tmp[5280]*kernel[0]+tmp[5281]*kernel[1]+tmp[5282]*kernel[2]+tmp[5380]*kernel[3]+tmp[5381]*kernel[4]+tmp[5382]*kernel[5]+tmp[5480]*kernel[6]+tmp[5481]*kernel[7]+tmp[5482]*kernel[8];
				ans[5382]<=tmp[5281]*kernel[0]+tmp[5282]*kernel[1]+tmp[5283]*kernel[2]+tmp[5381]*kernel[3]+tmp[5382]*kernel[4]+tmp[5383]*kernel[5]+tmp[5481]*kernel[6]+tmp[5482]*kernel[7]+tmp[5483]*kernel[8];
				ans[5383]<=tmp[5282]*kernel[0]+tmp[5283]*kernel[1]+tmp[5284]*kernel[2]+tmp[5382]*kernel[3]+tmp[5383]*kernel[4]+tmp[5384]*kernel[5]+tmp[5482]*kernel[6]+tmp[5483]*kernel[7]+tmp[5484]*kernel[8];
				ans[5384]<=tmp[5283]*kernel[0]+tmp[5284]*kernel[1]+tmp[5285]*kernel[2]+tmp[5383]*kernel[3]+tmp[5384]*kernel[4]+tmp[5385]*kernel[5]+tmp[5483]*kernel[6]+tmp[5484]*kernel[7]+tmp[5485]*kernel[8];
				ans[5385]<=tmp[5284]*kernel[0]+tmp[5285]*kernel[1]+tmp[5286]*kernel[2]+tmp[5384]*kernel[3]+tmp[5385]*kernel[4]+tmp[5386]*kernel[5]+tmp[5484]*kernel[6]+tmp[5485]*kernel[7]+tmp[5486]*kernel[8];
				ans[5386]<=tmp[5285]*kernel[0]+tmp[5286]*kernel[1]+tmp[5287]*kernel[2]+tmp[5385]*kernel[3]+tmp[5386]*kernel[4]+tmp[5387]*kernel[5]+tmp[5485]*kernel[6]+tmp[5486]*kernel[7]+tmp[5487]*kernel[8];
				ans[5387]<=tmp[5286]*kernel[0]+tmp[5287]*kernel[1]+tmp[5288]*kernel[2]+tmp[5386]*kernel[3]+tmp[5387]*kernel[4]+tmp[5388]*kernel[5]+tmp[5486]*kernel[6]+tmp[5487]*kernel[7]+tmp[5488]*kernel[8];
				ans[5388]<=tmp[5287]*kernel[0]+tmp[5288]*kernel[1]+tmp[5289]*kernel[2]+tmp[5387]*kernel[3]+tmp[5388]*kernel[4]+tmp[5389]*kernel[5]+tmp[5487]*kernel[6]+tmp[5488]*kernel[7]+tmp[5489]*kernel[8];
				ans[5389]<=tmp[5288]*kernel[0]+tmp[5289]*kernel[1]+tmp[5290]*kernel[2]+tmp[5388]*kernel[3]+tmp[5389]*kernel[4]+tmp[5390]*kernel[5]+tmp[5488]*kernel[6]+tmp[5489]*kernel[7]+tmp[5490]*kernel[8];
				ans[5390]<=tmp[5289]*kernel[0]+tmp[5290]*kernel[1]+tmp[5291]*kernel[2]+tmp[5389]*kernel[3]+tmp[5390]*kernel[4]+tmp[5391]*kernel[5]+tmp[5489]*kernel[6]+tmp[5490]*kernel[7]+tmp[5491]*kernel[8];
				ans[5391]<=tmp[5290]*kernel[0]+tmp[5291]*kernel[1]+tmp[5292]*kernel[2]+tmp[5390]*kernel[3]+tmp[5391]*kernel[4]+tmp[5392]*kernel[5]+tmp[5490]*kernel[6]+tmp[5491]*kernel[7]+tmp[5492]*kernel[8];
				ans[5392]<=tmp[5291]*kernel[0]+tmp[5292]*kernel[1]+tmp[5293]*kernel[2]+tmp[5391]*kernel[3]+tmp[5392]*kernel[4]+tmp[5393]*kernel[5]+tmp[5491]*kernel[6]+tmp[5492]*kernel[7]+tmp[5493]*kernel[8];
				ans[5393]<=tmp[5292]*kernel[0]+tmp[5293]*kernel[1]+tmp[5294]*kernel[2]+tmp[5392]*kernel[3]+tmp[5393]*kernel[4]+tmp[5394]*kernel[5]+tmp[5492]*kernel[6]+tmp[5493]*kernel[7]+tmp[5494]*kernel[8];
				ans[5394]<=tmp[5293]*kernel[0]+tmp[5294]*kernel[1]+tmp[5295]*kernel[2]+tmp[5393]*kernel[3]+tmp[5394]*kernel[4]+tmp[5395]*kernel[5]+tmp[5493]*kernel[6]+tmp[5494]*kernel[7]+tmp[5495]*kernel[8];
				ans[5395]<=tmp[5294]*kernel[0]+tmp[5295]*kernel[1]+tmp[5296]*kernel[2]+tmp[5394]*kernel[3]+tmp[5395]*kernel[4]+tmp[5396]*kernel[5]+tmp[5494]*kernel[6]+tmp[5495]*kernel[7]+tmp[5496]*kernel[8];
				ans[5396]<=tmp[5295]*kernel[0]+tmp[5296]*kernel[1]+tmp[5297]*kernel[2]+tmp[5395]*kernel[3]+tmp[5396]*kernel[4]+tmp[5397]*kernel[5]+tmp[5495]*kernel[6]+tmp[5496]*kernel[7]+tmp[5497]*kernel[8];
				ans[5397]<=tmp[5296]*kernel[0]+tmp[5297]*kernel[1]+tmp[5298]*kernel[2]+tmp[5396]*kernel[3]+tmp[5397]*kernel[4]+tmp[5398]*kernel[5]+tmp[5496]*kernel[6]+tmp[5497]*kernel[7]+tmp[5498]*kernel[8];
				ans[5398]<=tmp[5297]*kernel[0]+tmp[5298]*kernel[1]+tmp[5299]*kernel[2]+tmp[5397]*kernel[3]+tmp[5398]*kernel[4]+tmp[5399]*kernel[5]+tmp[5497]*kernel[6]+tmp[5498]*kernel[7]+tmp[5499]*kernel[8];
				ans[5399]<=tmp[5298]*kernel[0]+tmp[5299]*kernel[1]+tmp[5398]*kernel[3]+tmp[5399]*kernel[4]+tmp[5498]*kernel[6]+tmp[5499]*kernel[7];
				ans[5400]<=tmp[5300]*kernel[1]+tmp[5301]*kernel[2]+tmp[5400]*kernel[4]+tmp[5401]*kernel[5]+tmp[5500]*kernel[7]+tmp[5501]*kernel[8];
				ans[5401]<=tmp[5300]*kernel[0]+tmp[5301]*kernel[1]+tmp[5302]*kernel[2]+tmp[5400]*kernel[3]+tmp[5401]*kernel[4]+tmp[5402]*kernel[5]+tmp[5500]*kernel[6]+tmp[5501]*kernel[7]+tmp[5502]*kernel[8];
				ans[5402]<=tmp[5301]*kernel[0]+tmp[5302]*kernel[1]+tmp[5303]*kernel[2]+tmp[5401]*kernel[3]+tmp[5402]*kernel[4]+tmp[5403]*kernel[5]+tmp[5501]*kernel[6]+tmp[5502]*kernel[7]+tmp[5503]*kernel[8];
				ans[5403]<=tmp[5302]*kernel[0]+tmp[5303]*kernel[1]+tmp[5304]*kernel[2]+tmp[5402]*kernel[3]+tmp[5403]*kernel[4]+tmp[5404]*kernel[5]+tmp[5502]*kernel[6]+tmp[5503]*kernel[7]+tmp[5504]*kernel[8];
				ans[5404]<=tmp[5303]*kernel[0]+tmp[5304]*kernel[1]+tmp[5305]*kernel[2]+tmp[5403]*kernel[3]+tmp[5404]*kernel[4]+tmp[5405]*kernel[5]+tmp[5503]*kernel[6]+tmp[5504]*kernel[7]+tmp[5505]*kernel[8];
				ans[5405]<=tmp[5304]*kernel[0]+tmp[5305]*kernel[1]+tmp[5306]*kernel[2]+tmp[5404]*kernel[3]+tmp[5405]*kernel[4]+tmp[5406]*kernel[5]+tmp[5504]*kernel[6]+tmp[5505]*kernel[7]+tmp[5506]*kernel[8];
				ans[5406]<=tmp[5305]*kernel[0]+tmp[5306]*kernel[1]+tmp[5307]*kernel[2]+tmp[5405]*kernel[3]+tmp[5406]*kernel[4]+tmp[5407]*kernel[5]+tmp[5505]*kernel[6]+tmp[5506]*kernel[7]+tmp[5507]*kernel[8];
				ans[5407]<=tmp[5306]*kernel[0]+tmp[5307]*kernel[1]+tmp[5308]*kernel[2]+tmp[5406]*kernel[3]+tmp[5407]*kernel[4]+tmp[5408]*kernel[5]+tmp[5506]*kernel[6]+tmp[5507]*kernel[7]+tmp[5508]*kernel[8];
				ans[5408]<=tmp[5307]*kernel[0]+tmp[5308]*kernel[1]+tmp[5309]*kernel[2]+tmp[5407]*kernel[3]+tmp[5408]*kernel[4]+tmp[5409]*kernel[5]+tmp[5507]*kernel[6]+tmp[5508]*kernel[7]+tmp[5509]*kernel[8];
				ans[5409]<=tmp[5308]*kernel[0]+tmp[5309]*kernel[1]+tmp[5310]*kernel[2]+tmp[5408]*kernel[3]+tmp[5409]*kernel[4]+tmp[5410]*kernel[5]+tmp[5508]*kernel[6]+tmp[5509]*kernel[7]+tmp[5510]*kernel[8];
				ans[5410]<=tmp[5309]*kernel[0]+tmp[5310]*kernel[1]+tmp[5311]*kernel[2]+tmp[5409]*kernel[3]+tmp[5410]*kernel[4]+tmp[5411]*kernel[5]+tmp[5509]*kernel[6]+tmp[5510]*kernel[7]+tmp[5511]*kernel[8];
				ans[5411]<=tmp[5310]*kernel[0]+tmp[5311]*kernel[1]+tmp[5312]*kernel[2]+tmp[5410]*kernel[3]+tmp[5411]*kernel[4]+tmp[5412]*kernel[5]+tmp[5510]*kernel[6]+tmp[5511]*kernel[7]+tmp[5512]*kernel[8];
				ans[5412]<=tmp[5311]*kernel[0]+tmp[5312]*kernel[1]+tmp[5313]*kernel[2]+tmp[5411]*kernel[3]+tmp[5412]*kernel[4]+tmp[5413]*kernel[5]+tmp[5511]*kernel[6]+tmp[5512]*kernel[7]+tmp[5513]*kernel[8];
				ans[5413]<=tmp[5312]*kernel[0]+tmp[5313]*kernel[1]+tmp[5314]*kernel[2]+tmp[5412]*kernel[3]+tmp[5413]*kernel[4]+tmp[5414]*kernel[5]+tmp[5512]*kernel[6]+tmp[5513]*kernel[7]+tmp[5514]*kernel[8];
				ans[5414]<=tmp[5313]*kernel[0]+tmp[5314]*kernel[1]+tmp[5315]*kernel[2]+tmp[5413]*kernel[3]+tmp[5414]*kernel[4]+tmp[5415]*kernel[5]+tmp[5513]*kernel[6]+tmp[5514]*kernel[7]+tmp[5515]*kernel[8];
				ans[5415]<=tmp[5314]*kernel[0]+tmp[5315]*kernel[1]+tmp[5316]*kernel[2]+tmp[5414]*kernel[3]+tmp[5415]*kernel[4]+tmp[5416]*kernel[5]+tmp[5514]*kernel[6]+tmp[5515]*kernel[7]+tmp[5516]*kernel[8];
				ans[5416]<=tmp[5315]*kernel[0]+tmp[5316]*kernel[1]+tmp[5317]*kernel[2]+tmp[5415]*kernel[3]+tmp[5416]*kernel[4]+tmp[5417]*kernel[5]+tmp[5515]*kernel[6]+tmp[5516]*kernel[7]+tmp[5517]*kernel[8];
				ans[5417]<=tmp[5316]*kernel[0]+tmp[5317]*kernel[1]+tmp[5318]*kernel[2]+tmp[5416]*kernel[3]+tmp[5417]*kernel[4]+tmp[5418]*kernel[5]+tmp[5516]*kernel[6]+tmp[5517]*kernel[7]+tmp[5518]*kernel[8];
				ans[5418]<=tmp[5317]*kernel[0]+tmp[5318]*kernel[1]+tmp[5319]*kernel[2]+tmp[5417]*kernel[3]+tmp[5418]*kernel[4]+tmp[5419]*kernel[5]+tmp[5517]*kernel[6]+tmp[5518]*kernel[7]+tmp[5519]*kernel[8];
				ans[5419]<=tmp[5318]*kernel[0]+tmp[5319]*kernel[1]+tmp[5320]*kernel[2]+tmp[5418]*kernel[3]+tmp[5419]*kernel[4]+tmp[5420]*kernel[5]+tmp[5518]*kernel[6]+tmp[5519]*kernel[7]+tmp[5520]*kernel[8];
				ans[5420]<=tmp[5319]*kernel[0]+tmp[5320]*kernel[1]+tmp[5321]*kernel[2]+tmp[5419]*kernel[3]+tmp[5420]*kernel[4]+tmp[5421]*kernel[5]+tmp[5519]*kernel[6]+tmp[5520]*kernel[7]+tmp[5521]*kernel[8];
				ans[5421]<=tmp[5320]*kernel[0]+tmp[5321]*kernel[1]+tmp[5322]*kernel[2]+tmp[5420]*kernel[3]+tmp[5421]*kernel[4]+tmp[5422]*kernel[5]+tmp[5520]*kernel[6]+tmp[5521]*kernel[7]+tmp[5522]*kernel[8];
				ans[5422]<=tmp[5321]*kernel[0]+tmp[5322]*kernel[1]+tmp[5323]*kernel[2]+tmp[5421]*kernel[3]+tmp[5422]*kernel[4]+tmp[5423]*kernel[5]+tmp[5521]*kernel[6]+tmp[5522]*kernel[7]+tmp[5523]*kernel[8];
				ans[5423]<=tmp[5322]*kernel[0]+tmp[5323]*kernel[1]+tmp[5324]*kernel[2]+tmp[5422]*kernel[3]+tmp[5423]*kernel[4]+tmp[5424]*kernel[5]+tmp[5522]*kernel[6]+tmp[5523]*kernel[7]+tmp[5524]*kernel[8];
				ans[5424]<=tmp[5323]*kernel[0]+tmp[5324]*kernel[1]+tmp[5325]*kernel[2]+tmp[5423]*kernel[3]+tmp[5424]*kernel[4]+tmp[5425]*kernel[5]+tmp[5523]*kernel[6]+tmp[5524]*kernel[7]+tmp[5525]*kernel[8];
				ans[5425]<=tmp[5324]*kernel[0]+tmp[5325]*kernel[1]+tmp[5326]*kernel[2]+tmp[5424]*kernel[3]+tmp[5425]*kernel[4]+tmp[5426]*kernel[5]+tmp[5524]*kernel[6]+tmp[5525]*kernel[7]+tmp[5526]*kernel[8];
				ans[5426]<=tmp[5325]*kernel[0]+tmp[5326]*kernel[1]+tmp[5327]*kernel[2]+tmp[5425]*kernel[3]+tmp[5426]*kernel[4]+tmp[5427]*kernel[5]+tmp[5525]*kernel[6]+tmp[5526]*kernel[7]+tmp[5527]*kernel[8];
				ans[5427]<=tmp[5326]*kernel[0]+tmp[5327]*kernel[1]+tmp[5328]*kernel[2]+tmp[5426]*kernel[3]+tmp[5427]*kernel[4]+tmp[5428]*kernel[5]+tmp[5526]*kernel[6]+tmp[5527]*kernel[7]+tmp[5528]*kernel[8];
				ans[5428]<=tmp[5327]*kernel[0]+tmp[5328]*kernel[1]+tmp[5329]*kernel[2]+tmp[5427]*kernel[3]+tmp[5428]*kernel[4]+tmp[5429]*kernel[5]+tmp[5527]*kernel[6]+tmp[5528]*kernel[7]+tmp[5529]*kernel[8];
				ans[5429]<=tmp[5328]*kernel[0]+tmp[5329]*kernel[1]+tmp[5330]*kernel[2]+tmp[5428]*kernel[3]+tmp[5429]*kernel[4]+tmp[5430]*kernel[5]+tmp[5528]*kernel[6]+tmp[5529]*kernel[7]+tmp[5530]*kernel[8];
				ans[5430]<=tmp[5329]*kernel[0]+tmp[5330]*kernel[1]+tmp[5331]*kernel[2]+tmp[5429]*kernel[3]+tmp[5430]*kernel[4]+tmp[5431]*kernel[5]+tmp[5529]*kernel[6]+tmp[5530]*kernel[7]+tmp[5531]*kernel[8];
				ans[5431]<=tmp[5330]*kernel[0]+tmp[5331]*kernel[1]+tmp[5332]*kernel[2]+tmp[5430]*kernel[3]+tmp[5431]*kernel[4]+tmp[5432]*kernel[5]+tmp[5530]*kernel[6]+tmp[5531]*kernel[7]+tmp[5532]*kernel[8];
				ans[5432]<=tmp[5331]*kernel[0]+tmp[5332]*kernel[1]+tmp[5333]*kernel[2]+tmp[5431]*kernel[3]+tmp[5432]*kernel[4]+tmp[5433]*kernel[5]+tmp[5531]*kernel[6]+tmp[5532]*kernel[7]+tmp[5533]*kernel[8];
				ans[5433]<=tmp[5332]*kernel[0]+tmp[5333]*kernel[1]+tmp[5334]*kernel[2]+tmp[5432]*kernel[3]+tmp[5433]*kernel[4]+tmp[5434]*kernel[5]+tmp[5532]*kernel[6]+tmp[5533]*kernel[7]+tmp[5534]*kernel[8];
				ans[5434]<=tmp[5333]*kernel[0]+tmp[5334]*kernel[1]+tmp[5335]*kernel[2]+tmp[5433]*kernel[3]+tmp[5434]*kernel[4]+tmp[5435]*kernel[5]+tmp[5533]*kernel[6]+tmp[5534]*kernel[7]+tmp[5535]*kernel[8];
				ans[5435]<=tmp[5334]*kernel[0]+tmp[5335]*kernel[1]+tmp[5336]*kernel[2]+tmp[5434]*kernel[3]+tmp[5435]*kernel[4]+tmp[5436]*kernel[5]+tmp[5534]*kernel[6]+tmp[5535]*kernel[7]+tmp[5536]*kernel[8];
				ans[5436]<=tmp[5335]*kernel[0]+tmp[5336]*kernel[1]+tmp[5337]*kernel[2]+tmp[5435]*kernel[3]+tmp[5436]*kernel[4]+tmp[5437]*kernel[5]+tmp[5535]*kernel[6]+tmp[5536]*kernel[7]+tmp[5537]*kernel[8];
				ans[5437]<=tmp[5336]*kernel[0]+tmp[5337]*kernel[1]+tmp[5338]*kernel[2]+tmp[5436]*kernel[3]+tmp[5437]*kernel[4]+tmp[5438]*kernel[5]+tmp[5536]*kernel[6]+tmp[5537]*kernel[7]+tmp[5538]*kernel[8];
				ans[5438]<=tmp[5337]*kernel[0]+tmp[5338]*kernel[1]+tmp[5339]*kernel[2]+tmp[5437]*kernel[3]+tmp[5438]*kernel[4]+tmp[5439]*kernel[5]+tmp[5537]*kernel[6]+tmp[5538]*kernel[7]+tmp[5539]*kernel[8];
				ans[5439]<=tmp[5338]*kernel[0]+tmp[5339]*kernel[1]+tmp[5340]*kernel[2]+tmp[5438]*kernel[3]+tmp[5439]*kernel[4]+tmp[5440]*kernel[5]+tmp[5538]*kernel[6]+tmp[5539]*kernel[7]+tmp[5540]*kernel[8];
				ans[5440]<=tmp[5339]*kernel[0]+tmp[5340]*kernel[1]+tmp[5341]*kernel[2]+tmp[5439]*kernel[3]+tmp[5440]*kernel[4]+tmp[5441]*kernel[5]+tmp[5539]*kernel[6]+tmp[5540]*kernel[7]+tmp[5541]*kernel[8];
				ans[5441]<=tmp[5340]*kernel[0]+tmp[5341]*kernel[1]+tmp[5342]*kernel[2]+tmp[5440]*kernel[3]+tmp[5441]*kernel[4]+tmp[5442]*kernel[5]+tmp[5540]*kernel[6]+tmp[5541]*kernel[7]+tmp[5542]*kernel[8];
				ans[5442]<=tmp[5341]*kernel[0]+tmp[5342]*kernel[1]+tmp[5343]*kernel[2]+tmp[5441]*kernel[3]+tmp[5442]*kernel[4]+tmp[5443]*kernel[5]+tmp[5541]*kernel[6]+tmp[5542]*kernel[7]+tmp[5543]*kernel[8];
				ans[5443]<=tmp[5342]*kernel[0]+tmp[5343]*kernel[1]+tmp[5344]*kernel[2]+tmp[5442]*kernel[3]+tmp[5443]*kernel[4]+tmp[5444]*kernel[5]+tmp[5542]*kernel[6]+tmp[5543]*kernel[7]+tmp[5544]*kernel[8];
				ans[5444]<=tmp[5343]*kernel[0]+tmp[5344]*kernel[1]+tmp[5345]*kernel[2]+tmp[5443]*kernel[3]+tmp[5444]*kernel[4]+tmp[5445]*kernel[5]+tmp[5543]*kernel[6]+tmp[5544]*kernel[7]+tmp[5545]*kernel[8];
				ans[5445]<=tmp[5344]*kernel[0]+tmp[5345]*kernel[1]+tmp[5346]*kernel[2]+tmp[5444]*kernel[3]+tmp[5445]*kernel[4]+tmp[5446]*kernel[5]+tmp[5544]*kernel[6]+tmp[5545]*kernel[7]+tmp[5546]*kernel[8];
				ans[5446]<=tmp[5345]*kernel[0]+tmp[5346]*kernel[1]+tmp[5347]*kernel[2]+tmp[5445]*kernel[3]+tmp[5446]*kernel[4]+tmp[5447]*kernel[5]+tmp[5545]*kernel[6]+tmp[5546]*kernel[7]+tmp[5547]*kernel[8];
				ans[5447]<=tmp[5346]*kernel[0]+tmp[5347]*kernel[1]+tmp[5348]*kernel[2]+tmp[5446]*kernel[3]+tmp[5447]*kernel[4]+tmp[5448]*kernel[5]+tmp[5546]*kernel[6]+tmp[5547]*kernel[7]+tmp[5548]*kernel[8];
				ans[5448]<=tmp[5347]*kernel[0]+tmp[5348]*kernel[1]+tmp[5349]*kernel[2]+tmp[5447]*kernel[3]+tmp[5448]*kernel[4]+tmp[5449]*kernel[5]+tmp[5547]*kernel[6]+tmp[5548]*kernel[7]+tmp[5549]*kernel[8];
				ans[5449]<=tmp[5348]*kernel[0]+tmp[5349]*kernel[1]+tmp[5350]*kernel[2]+tmp[5448]*kernel[3]+tmp[5449]*kernel[4]+tmp[5450]*kernel[5]+tmp[5548]*kernel[6]+tmp[5549]*kernel[7]+tmp[5550]*kernel[8];
				ans[5450]<=tmp[5349]*kernel[0]+tmp[5350]*kernel[1]+tmp[5351]*kernel[2]+tmp[5449]*kernel[3]+tmp[5450]*kernel[4]+tmp[5451]*kernel[5]+tmp[5549]*kernel[6]+tmp[5550]*kernel[7]+tmp[5551]*kernel[8];
				ans[5451]<=tmp[5350]*kernel[0]+tmp[5351]*kernel[1]+tmp[5352]*kernel[2]+tmp[5450]*kernel[3]+tmp[5451]*kernel[4]+tmp[5452]*kernel[5]+tmp[5550]*kernel[6]+tmp[5551]*kernel[7]+tmp[5552]*kernel[8];
				ans[5452]<=tmp[5351]*kernel[0]+tmp[5352]*kernel[1]+tmp[5353]*kernel[2]+tmp[5451]*kernel[3]+tmp[5452]*kernel[4]+tmp[5453]*kernel[5]+tmp[5551]*kernel[6]+tmp[5552]*kernel[7]+tmp[5553]*kernel[8];
				ans[5453]<=tmp[5352]*kernel[0]+tmp[5353]*kernel[1]+tmp[5354]*kernel[2]+tmp[5452]*kernel[3]+tmp[5453]*kernel[4]+tmp[5454]*kernel[5]+tmp[5552]*kernel[6]+tmp[5553]*kernel[7]+tmp[5554]*kernel[8];
				ans[5454]<=tmp[5353]*kernel[0]+tmp[5354]*kernel[1]+tmp[5355]*kernel[2]+tmp[5453]*kernel[3]+tmp[5454]*kernel[4]+tmp[5455]*kernel[5]+tmp[5553]*kernel[6]+tmp[5554]*kernel[7]+tmp[5555]*kernel[8];
				ans[5455]<=tmp[5354]*kernel[0]+tmp[5355]*kernel[1]+tmp[5356]*kernel[2]+tmp[5454]*kernel[3]+tmp[5455]*kernel[4]+tmp[5456]*kernel[5]+tmp[5554]*kernel[6]+tmp[5555]*kernel[7]+tmp[5556]*kernel[8];
				ans[5456]<=tmp[5355]*kernel[0]+tmp[5356]*kernel[1]+tmp[5357]*kernel[2]+tmp[5455]*kernel[3]+tmp[5456]*kernel[4]+tmp[5457]*kernel[5]+tmp[5555]*kernel[6]+tmp[5556]*kernel[7]+tmp[5557]*kernel[8];
				ans[5457]<=tmp[5356]*kernel[0]+tmp[5357]*kernel[1]+tmp[5358]*kernel[2]+tmp[5456]*kernel[3]+tmp[5457]*kernel[4]+tmp[5458]*kernel[5]+tmp[5556]*kernel[6]+tmp[5557]*kernel[7]+tmp[5558]*kernel[8];
				ans[5458]<=tmp[5357]*kernel[0]+tmp[5358]*kernel[1]+tmp[5359]*kernel[2]+tmp[5457]*kernel[3]+tmp[5458]*kernel[4]+tmp[5459]*kernel[5]+tmp[5557]*kernel[6]+tmp[5558]*kernel[7]+tmp[5559]*kernel[8];
				ans[5459]<=tmp[5358]*kernel[0]+tmp[5359]*kernel[1]+tmp[5360]*kernel[2]+tmp[5458]*kernel[3]+tmp[5459]*kernel[4]+tmp[5460]*kernel[5]+tmp[5558]*kernel[6]+tmp[5559]*kernel[7]+tmp[5560]*kernel[8];
				ans[5460]<=tmp[5359]*kernel[0]+tmp[5360]*kernel[1]+tmp[5361]*kernel[2]+tmp[5459]*kernel[3]+tmp[5460]*kernel[4]+tmp[5461]*kernel[5]+tmp[5559]*kernel[6]+tmp[5560]*kernel[7]+tmp[5561]*kernel[8];
				ans[5461]<=tmp[5360]*kernel[0]+tmp[5361]*kernel[1]+tmp[5362]*kernel[2]+tmp[5460]*kernel[3]+tmp[5461]*kernel[4]+tmp[5462]*kernel[5]+tmp[5560]*kernel[6]+tmp[5561]*kernel[7]+tmp[5562]*kernel[8];
				ans[5462]<=tmp[5361]*kernel[0]+tmp[5362]*kernel[1]+tmp[5363]*kernel[2]+tmp[5461]*kernel[3]+tmp[5462]*kernel[4]+tmp[5463]*kernel[5]+tmp[5561]*kernel[6]+tmp[5562]*kernel[7]+tmp[5563]*kernel[8];
				ans[5463]<=tmp[5362]*kernel[0]+tmp[5363]*kernel[1]+tmp[5364]*kernel[2]+tmp[5462]*kernel[3]+tmp[5463]*kernel[4]+tmp[5464]*kernel[5]+tmp[5562]*kernel[6]+tmp[5563]*kernel[7]+tmp[5564]*kernel[8];
				ans[5464]<=tmp[5363]*kernel[0]+tmp[5364]*kernel[1]+tmp[5365]*kernel[2]+tmp[5463]*kernel[3]+tmp[5464]*kernel[4]+tmp[5465]*kernel[5]+tmp[5563]*kernel[6]+tmp[5564]*kernel[7]+tmp[5565]*kernel[8];
				ans[5465]<=tmp[5364]*kernel[0]+tmp[5365]*kernel[1]+tmp[5366]*kernel[2]+tmp[5464]*kernel[3]+tmp[5465]*kernel[4]+tmp[5466]*kernel[5]+tmp[5564]*kernel[6]+tmp[5565]*kernel[7]+tmp[5566]*kernel[8];
				ans[5466]<=tmp[5365]*kernel[0]+tmp[5366]*kernel[1]+tmp[5367]*kernel[2]+tmp[5465]*kernel[3]+tmp[5466]*kernel[4]+tmp[5467]*kernel[5]+tmp[5565]*kernel[6]+tmp[5566]*kernel[7]+tmp[5567]*kernel[8];
				ans[5467]<=tmp[5366]*kernel[0]+tmp[5367]*kernel[1]+tmp[5368]*kernel[2]+tmp[5466]*kernel[3]+tmp[5467]*kernel[4]+tmp[5468]*kernel[5]+tmp[5566]*kernel[6]+tmp[5567]*kernel[7]+tmp[5568]*kernel[8];
				ans[5468]<=tmp[5367]*kernel[0]+tmp[5368]*kernel[1]+tmp[5369]*kernel[2]+tmp[5467]*kernel[3]+tmp[5468]*kernel[4]+tmp[5469]*kernel[5]+tmp[5567]*kernel[6]+tmp[5568]*kernel[7]+tmp[5569]*kernel[8];
				ans[5469]<=tmp[5368]*kernel[0]+tmp[5369]*kernel[1]+tmp[5370]*kernel[2]+tmp[5468]*kernel[3]+tmp[5469]*kernel[4]+tmp[5470]*kernel[5]+tmp[5568]*kernel[6]+tmp[5569]*kernel[7]+tmp[5570]*kernel[8];
				ans[5470]<=tmp[5369]*kernel[0]+tmp[5370]*kernel[1]+tmp[5371]*kernel[2]+tmp[5469]*kernel[3]+tmp[5470]*kernel[4]+tmp[5471]*kernel[5]+tmp[5569]*kernel[6]+tmp[5570]*kernel[7]+tmp[5571]*kernel[8];
				ans[5471]<=tmp[5370]*kernel[0]+tmp[5371]*kernel[1]+tmp[5372]*kernel[2]+tmp[5470]*kernel[3]+tmp[5471]*kernel[4]+tmp[5472]*kernel[5]+tmp[5570]*kernel[6]+tmp[5571]*kernel[7]+tmp[5572]*kernel[8];
				ans[5472]<=tmp[5371]*kernel[0]+tmp[5372]*kernel[1]+tmp[5373]*kernel[2]+tmp[5471]*kernel[3]+tmp[5472]*kernel[4]+tmp[5473]*kernel[5]+tmp[5571]*kernel[6]+tmp[5572]*kernel[7]+tmp[5573]*kernel[8];
				ans[5473]<=tmp[5372]*kernel[0]+tmp[5373]*kernel[1]+tmp[5374]*kernel[2]+tmp[5472]*kernel[3]+tmp[5473]*kernel[4]+tmp[5474]*kernel[5]+tmp[5572]*kernel[6]+tmp[5573]*kernel[7]+tmp[5574]*kernel[8];
				ans[5474]<=tmp[5373]*kernel[0]+tmp[5374]*kernel[1]+tmp[5375]*kernel[2]+tmp[5473]*kernel[3]+tmp[5474]*kernel[4]+tmp[5475]*kernel[5]+tmp[5573]*kernel[6]+tmp[5574]*kernel[7]+tmp[5575]*kernel[8];
				ans[5475]<=tmp[5374]*kernel[0]+tmp[5375]*kernel[1]+tmp[5376]*kernel[2]+tmp[5474]*kernel[3]+tmp[5475]*kernel[4]+tmp[5476]*kernel[5]+tmp[5574]*kernel[6]+tmp[5575]*kernel[7]+tmp[5576]*kernel[8];
				ans[5476]<=tmp[5375]*kernel[0]+tmp[5376]*kernel[1]+tmp[5377]*kernel[2]+tmp[5475]*kernel[3]+tmp[5476]*kernel[4]+tmp[5477]*kernel[5]+tmp[5575]*kernel[6]+tmp[5576]*kernel[7]+tmp[5577]*kernel[8];
				ans[5477]<=tmp[5376]*kernel[0]+tmp[5377]*kernel[1]+tmp[5378]*kernel[2]+tmp[5476]*kernel[3]+tmp[5477]*kernel[4]+tmp[5478]*kernel[5]+tmp[5576]*kernel[6]+tmp[5577]*kernel[7]+tmp[5578]*kernel[8];
				ans[5478]<=tmp[5377]*kernel[0]+tmp[5378]*kernel[1]+tmp[5379]*kernel[2]+tmp[5477]*kernel[3]+tmp[5478]*kernel[4]+tmp[5479]*kernel[5]+tmp[5577]*kernel[6]+tmp[5578]*kernel[7]+tmp[5579]*kernel[8];
				ans[5479]<=tmp[5378]*kernel[0]+tmp[5379]*kernel[1]+tmp[5380]*kernel[2]+tmp[5478]*kernel[3]+tmp[5479]*kernel[4]+tmp[5480]*kernel[5]+tmp[5578]*kernel[6]+tmp[5579]*kernel[7]+tmp[5580]*kernel[8];
				ans[5480]<=tmp[5379]*kernel[0]+tmp[5380]*kernel[1]+tmp[5381]*kernel[2]+tmp[5479]*kernel[3]+tmp[5480]*kernel[4]+tmp[5481]*kernel[5]+tmp[5579]*kernel[6]+tmp[5580]*kernel[7]+tmp[5581]*kernel[8];
				ans[5481]<=tmp[5380]*kernel[0]+tmp[5381]*kernel[1]+tmp[5382]*kernel[2]+tmp[5480]*kernel[3]+tmp[5481]*kernel[4]+tmp[5482]*kernel[5]+tmp[5580]*kernel[6]+tmp[5581]*kernel[7]+tmp[5582]*kernel[8];
				ans[5482]<=tmp[5381]*kernel[0]+tmp[5382]*kernel[1]+tmp[5383]*kernel[2]+tmp[5481]*kernel[3]+tmp[5482]*kernel[4]+tmp[5483]*kernel[5]+tmp[5581]*kernel[6]+tmp[5582]*kernel[7]+tmp[5583]*kernel[8];
				ans[5483]<=tmp[5382]*kernel[0]+tmp[5383]*kernel[1]+tmp[5384]*kernel[2]+tmp[5482]*kernel[3]+tmp[5483]*kernel[4]+tmp[5484]*kernel[5]+tmp[5582]*kernel[6]+tmp[5583]*kernel[7]+tmp[5584]*kernel[8];
				ans[5484]<=tmp[5383]*kernel[0]+tmp[5384]*kernel[1]+tmp[5385]*kernel[2]+tmp[5483]*kernel[3]+tmp[5484]*kernel[4]+tmp[5485]*kernel[5]+tmp[5583]*kernel[6]+tmp[5584]*kernel[7]+tmp[5585]*kernel[8];
				ans[5485]<=tmp[5384]*kernel[0]+tmp[5385]*kernel[1]+tmp[5386]*kernel[2]+tmp[5484]*kernel[3]+tmp[5485]*kernel[4]+tmp[5486]*kernel[5]+tmp[5584]*kernel[6]+tmp[5585]*kernel[7]+tmp[5586]*kernel[8];
				ans[5486]<=tmp[5385]*kernel[0]+tmp[5386]*kernel[1]+tmp[5387]*kernel[2]+tmp[5485]*kernel[3]+tmp[5486]*kernel[4]+tmp[5487]*kernel[5]+tmp[5585]*kernel[6]+tmp[5586]*kernel[7]+tmp[5587]*kernel[8];
				ans[5487]<=tmp[5386]*kernel[0]+tmp[5387]*kernel[1]+tmp[5388]*kernel[2]+tmp[5486]*kernel[3]+tmp[5487]*kernel[4]+tmp[5488]*kernel[5]+tmp[5586]*kernel[6]+tmp[5587]*kernel[7]+tmp[5588]*kernel[8];
				ans[5488]<=tmp[5387]*kernel[0]+tmp[5388]*kernel[1]+tmp[5389]*kernel[2]+tmp[5487]*kernel[3]+tmp[5488]*kernel[4]+tmp[5489]*kernel[5]+tmp[5587]*kernel[6]+tmp[5588]*kernel[7]+tmp[5589]*kernel[8];
				ans[5489]<=tmp[5388]*kernel[0]+tmp[5389]*kernel[1]+tmp[5390]*kernel[2]+tmp[5488]*kernel[3]+tmp[5489]*kernel[4]+tmp[5490]*kernel[5]+tmp[5588]*kernel[6]+tmp[5589]*kernel[7]+tmp[5590]*kernel[8];
				ans[5490]<=tmp[5389]*kernel[0]+tmp[5390]*kernel[1]+tmp[5391]*kernel[2]+tmp[5489]*kernel[3]+tmp[5490]*kernel[4]+tmp[5491]*kernel[5]+tmp[5589]*kernel[6]+tmp[5590]*kernel[7]+tmp[5591]*kernel[8];
				ans[5491]<=tmp[5390]*kernel[0]+tmp[5391]*kernel[1]+tmp[5392]*kernel[2]+tmp[5490]*kernel[3]+tmp[5491]*kernel[4]+tmp[5492]*kernel[5]+tmp[5590]*kernel[6]+tmp[5591]*kernel[7]+tmp[5592]*kernel[8];
				ans[5492]<=tmp[5391]*kernel[0]+tmp[5392]*kernel[1]+tmp[5393]*kernel[2]+tmp[5491]*kernel[3]+tmp[5492]*kernel[4]+tmp[5493]*kernel[5]+tmp[5591]*kernel[6]+tmp[5592]*kernel[7]+tmp[5593]*kernel[8];
				ans[5493]<=tmp[5392]*kernel[0]+tmp[5393]*kernel[1]+tmp[5394]*kernel[2]+tmp[5492]*kernel[3]+tmp[5493]*kernel[4]+tmp[5494]*kernel[5]+tmp[5592]*kernel[6]+tmp[5593]*kernel[7]+tmp[5594]*kernel[8];
				ans[5494]<=tmp[5393]*kernel[0]+tmp[5394]*kernel[1]+tmp[5395]*kernel[2]+tmp[5493]*kernel[3]+tmp[5494]*kernel[4]+tmp[5495]*kernel[5]+tmp[5593]*kernel[6]+tmp[5594]*kernel[7]+tmp[5595]*kernel[8];
				ans[5495]<=tmp[5394]*kernel[0]+tmp[5395]*kernel[1]+tmp[5396]*kernel[2]+tmp[5494]*kernel[3]+tmp[5495]*kernel[4]+tmp[5496]*kernel[5]+tmp[5594]*kernel[6]+tmp[5595]*kernel[7]+tmp[5596]*kernel[8];
				ans[5496]<=tmp[5395]*kernel[0]+tmp[5396]*kernel[1]+tmp[5397]*kernel[2]+tmp[5495]*kernel[3]+tmp[5496]*kernel[4]+tmp[5497]*kernel[5]+tmp[5595]*kernel[6]+tmp[5596]*kernel[7]+tmp[5597]*kernel[8];
				ans[5497]<=tmp[5396]*kernel[0]+tmp[5397]*kernel[1]+tmp[5398]*kernel[2]+tmp[5496]*kernel[3]+tmp[5497]*kernel[4]+tmp[5498]*kernel[5]+tmp[5596]*kernel[6]+tmp[5597]*kernel[7]+tmp[5598]*kernel[8];
				ans[5498]<=tmp[5397]*kernel[0]+tmp[5398]*kernel[1]+tmp[5399]*kernel[2]+tmp[5497]*kernel[3]+tmp[5498]*kernel[4]+tmp[5499]*kernel[5]+tmp[5597]*kernel[6]+tmp[5598]*kernel[7]+tmp[5599]*kernel[8];
				ans[5499]<=tmp[5398]*kernel[0]+tmp[5399]*kernel[1]+tmp[5498]*kernel[3]+tmp[5499]*kernel[4]+tmp[5598]*kernel[6]+tmp[5599]*kernel[7];
				ans[5500]<=tmp[5400]*kernel[1]+tmp[5401]*kernel[2]+tmp[5500]*kernel[4]+tmp[5501]*kernel[5]+tmp[5600]*kernel[7]+tmp[5601]*kernel[8];
				ans[5501]<=tmp[5400]*kernel[0]+tmp[5401]*kernel[1]+tmp[5402]*kernel[2]+tmp[5500]*kernel[3]+tmp[5501]*kernel[4]+tmp[5502]*kernel[5]+tmp[5600]*kernel[6]+tmp[5601]*kernel[7]+tmp[5602]*kernel[8];
				ans[5502]<=tmp[5401]*kernel[0]+tmp[5402]*kernel[1]+tmp[5403]*kernel[2]+tmp[5501]*kernel[3]+tmp[5502]*kernel[4]+tmp[5503]*kernel[5]+tmp[5601]*kernel[6]+tmp[5602]*kernel[7]+tmp[5603]*kernel[8];
				ans[5503]<=tmp[5402]*kernel[0]+tmp[5403]*kernel[1]+tmp[5404]*kernel[2]+tmp[5502]*kernel[3]+tmp[5503]*kernel[4]+tmp[5504]*kernel[5]+tmp[5602]*kernel[6]+tmp[5603]*kernel[7]+tmp[5604]*kernel[8];
				ans[5504]<=tmp[5403]*kernel[0]+tmp[5404]*kernel[1]+tmp[5405]*kernel[2]+tmp[5503]*kernel[3]+tmp[5504]*kernel[4]+tmp[5505]*kernel[5]+tmp[5603]*kernel[6]+tmp[5604]*kernel[7]+tmp[5605]*kernel[8];
				ans[5505]<=tmp[5404]*kernel[0]+tmp[5405]*kernel[1]+tmp[5406]*kernel[2]+tmp[5504]*kernel[3]+tmp[5505]*kernel[4]+tmp[5506]*kernel[5]+tmp[5604]*kernel[6]+tmp[5605]*kernel[7]+tmp[5606]*kernel[8];
				ans[5506]<=tmp[5405]*kernel[0]+tmp[5406]*kernel[1]+tmp[5407]*kernel[2]+tmp[5505]*kernel[3]+tmp[5506]*kernel[4]+tmp[5507]*kernel[5]+tmp[5605]*kernel[6]+tmp[5606]*kernel[7]+tmp[5607]*kernel[8];
				ans[5507]<=tmp[5406]*kernel[0]+tmp[5407]*kernel[1]+tmp[5408]*kernel[2]+tmp[5506]*kernel[3]+tmp[5507]*kernel[4]+tmp[5508]*kernel[5]+tmp[5606]*kernel[6]+tmp[5607]*kernel[7]+tmp[5608]*kernel[8];
				ans[5508]<=tmp[5407]*kernel[0]+tmp[5408]*kernel[1]+tmp[5409]*kernel[2]+tmp[5507]*kernel[3]+tmp[5508]*kernel[4]+tmp[5509]*kernel[5]+tmp[5607]*kernel[6]+tmp[5608]*kernel[7]+tmp[5609]*kernel[8];
				ans[5509]<=tmp[5408]*kernel[0]+tmp[5409]*kernel[1]+tmp[5410]*kernel[2]+tmp[5508]*kernel[3]+tmp[5509]*kernel[4]+tmp[5510]*kernel[5]+tmp[5608]*kernel[6]+tmp[5609]*kernel[7]+tmp[5610]*kernel[8];
				ans[5510]<=tmp[5409]*kernel[0]+tmp[5410]*kernel[1]+tmp[5411]*kernel[2]+tmp[5509]*kernel[3]+tmp[5510]*kernel[4]+tmp[5511]*kernel[5]+tmp[5609]*kernel[6]+tmp[5610]*kernel[7]+tmp[5611]*kernel[8];
				ans[5511]<=tmp[5410]*kernel[0]+tmp[5411]*kernel[1]+tmp[5412]*kernel[2]+tmp[5510]*kernel[3]+tmp[5511]*kernel[4]+tmp[5512]*kernel[5]+tmp[5610]*kernel[6]+tmp[5611]*kernel[7]+tmp[5612]*kernel[8];
				ans[5512]<=tmp[5411]*kernel[0]+tmp[5412]*kernel[1]+tmp[5413]*kernel[2]+tmp[5511]*kernel[3]+tmp[5512]*kernel[4]+tmp[5513]*kernel[5]+tmp[5611]*kernel[6]+tmp[5612]*kernel[7]+tmp[5613]*kernel[8];
				ans[5513]<=tmp[5412]*kernel[0]+tmp[5413]*kernel[1]+tmp[5414]*kernel[2]+tmp[5512]*kernel[3]+tmp[5513]*kernel[4]+tmp[5514]*kernel[5]+tmp[5612]*kernel[6]+tmp[5613]*kernel[7]+tmp[5614]*kernel[8];
				ans[5514]<=tmp[5413]*kernel[0]+tmp[5414]*kernel[1]+tmp[5415]*kernel[2]+tmp[5513]*kernel[3]+tmp[5514]*kernel[4]+tmp[5515]*kernel[5]+tmp[5613]*kernel[6]+tmp[5614]*kernel[7]+tmp[5615]*kernel[8];
				ans[5515]<=tmp[5414]*kernel[0]+tmp[5415]*kernel[1]+tmp[5416]*kernel[2]+tmp[5514]*kernel[3]+tmp[5515]*kernel[4]+tmp[5516]*kernel[5]+tmp[5614]*kernel[6]+tmp[5615]*kernel[7]+tmp[5616]*kernel[8];
				ans[5516]<=tmp[5415]*kernel[0]+tmp[5416]*kernel[1]+tmp[5417]*kernel[2]+tmp[5515]*kernel[3]+tmp[5516]*kernel[4]+tmp[5517]*kernel[5]+tmp[5615]*kernel[6]+tmp[5616]*kernel[7]+tmp[5617]*kernel[8];
				ans[5517]<=tmp[5416]*kernel[0]+tmp[5417]*kernel[1]+tmp[5418]*kernel[2]+tmp[5516]*kernel[3]+tmp[5517]*kernel[4]+tmp[5518]*kernel[5]+tmp[5616]*kernel[6]+tmp[5617]*kernel[7]+tmp[5618]*kernel[8];
				ans[5518]<=tmp[5417]*kernel[0]+tmp[5418]*kernel[1]+tmp[5419]*kernel[2]+tmp[5517]*kernel[3]+tmp[5518]*kernel[4]+tmp[5519]*kernel[5]+tmp[5617]*kernel[6]+tmp[5618]*kernel[7]+tmp[5619]*kernel[8];
				ans[5519]<=tmp[5418]*kernel[0]+tmp[5419]*kernel[1]+tmp[5420]*kernel[2]+tmp[5518]*kernel[3]+tmp[5519]*kernel[4]+tmp[5520]*kernel[5]+tmp[5618]*kernel[6]+tmp[5619]*kernel[7]+tmp[5620]*kernel[8];
				ans[5520]<=tmp[5419]*kernel[0]+tmp[5420]*kernel[1]+tmp[5421]*kernel[2]+tmp[5519]*kernel[3]+tmp[5520]*kernel[4]+tmp[5521]*kernel[5]+tmp[5619]*kernel[6]+tmp[5620]*kernel[7]+tmp[5621]*kernel[8];
				ans[5521]<=tmp[5420]*kernel[0]+tmp[5421]*kernel[1]+tmp[5422]*kernel[2]+tmp[5520]*kernel[3]+tmp[5521]*kernel[4]+tmp[5522]*kernel[5]+tmp[5620]*kernel[6]+tmp[5621]*kernel[7]+tmp[5622]*kernel[8];
				ans[5522]<=tmp[5421]*kernel[0]+tmp[5422]*kernel[1]+tmp[5423]*kernel[2]+tmp[5521]*kernel[3]+tmp[5522]*kernel[4]+tmp[5523]*kernel[5]+tmp[5621]*kernel[6]+tmp[5622]*kernel[7]+tmp[5623]*kernel[8];
				ans[5523]<=tmp[5422]*kernel[0]+tmp[5423]*kernel[1]+tmp[5424]*kernel[2]+tmp[5522]*kernel[3]+tmp[5523]*kernel[4]+tmp[5524]*kernel[5]+tmp[5622]*kernel[6]+tmp[5623]*kernel[7]+tmp[5624]*kernel[8];
				ans[5524]<=tmp[5423]*kernel[0]+tmp[5424]*kernel[1]+tmp[5425]*kernel[2]+tmp[5523]*kernel[3]+tmp[5524]*kernel[4]+tmp[5525]*kernel[5]+tmp[5623]*kernel[6]+tmp[5624]*kernel[7]+tmp[5625]*kernel[8];
				ans[5525]<=tmp[5424]*kernel[0]+tmp[5425]*kernel[1]+tmp[5426]*kernel[2]+tmp[5524]*kernel[3]+tmp[5525]*kernel[4]+tmp[5526]*kernel[5]+tmp[5624]*kernel[6]+tmp[5625]*kernel[7]+tmp[5626]*kernel[8];
				ans[5526]<=tmp[5425]*kernel[0]+tmp[5426]*kernel[1]+tmp[5427]*kernel[2]+tmp[5525]*kernel[3]+tmp[5526]*kernel[4]+tmp[5527]*kernel[5]+tmp[5625]*kernel[6]+tmp[5626]*kernel[7]+tmp[5627]*kernel[8];
				ans[5527]<=tmp[5426]*kernel[0]+tmp[5427]*kernel[1]+tmp[5428]*kernel[2]+tmp[5526]*kernel[3]+tmp[5527]*kernel[4]+tmp[5528]*kernel[5]+tmp[5626]*kernel[6]+tmp[5627]*kernel[7]+tmp[5628]*kernel[8];
				ans[5528]<=tmp[5427]*kernel[0]+tmp[5428]*kernel[1]+tmp[5429]*kernel[2]+tmp[5527]*kernel[3]+tmp[5528]*kernel[4]+tmp[5529]*kernel[5]+tmp[5627]*kernel[6]+tmp[5628]*kernel[7]+tmp[5629]*kernel[8];
				ans[5529]<=tmp[5428]*kernel[0]+tmp[5429]*kernel[1]+tmp[5430]*kernel[2]+tmp[5528]*kernel[3]+tmp[5529]*kernel[4]+tmp[5530]*kernel[5]+tmp[5628]*kernel[6]+tmp[5629]*kernel[7]+tmp[5630]*kernel[8];
				ans[5530]<=tmp[5429]*kernel[0]+tmp[5430]*kernel[1]+tmp[5431]*kernel[2]+tmp[5529]*kernel[3]+tmp[5530]*kernel[4]+tmp[5531]*kernel[5]+tmp[5629]*kernel[6]+tmp[5630]*kernel[7]+tmp[5631]*kernel[8];
				ans[5531]<=tmp[5430]*kernel[0]+tmp[5431]*kernel[1]+tmp[5432]*kernel[2]+tmp[5530]*kernel[3]+tmp[5531]*kernel[4]+tmp[5532]*kernel[5]+tmp[5630]*kernel[6]+tmp[5631]*kernel[7]+tmp[5632]*kernel[8];
				ans[5532]<=tmp[5431]*kernel[0]+tmp[5432]*kernel[1]+tmp[5433]*kernel[2]+tmp[5531]*kernel[3]+tmp[5532]*kernel[4]+tmp[5533]*kernel[5]+tmp[5631]*kernel[6]+tmp[5632]*kernel[7]+tmp[5633]*kernel[8];
				ans[5533]<=tmp[5432]*kernel[0]+tmp[5433]*kernel[1]+tmp[5434]*kernel[2]+tmp[5532]*kernel[3]+tmp[5533]*kernel[4]+tmp[5534]*kernel[5]+tmp[5632]*kernel[6]+tmp[5633]*kernel[7]+tmp[5634]*kernel[8];
				ans[5534]<=tmp[5433]*kernel[0]+tmp[5434]*kernel[1]+tmp[5435]*kernel[2]+tmp[5533]*kernel[3]+tmp[5534]*kernel[4]+tmp[5535]*kernel[5]+tmp[5633]*kernel[6]+tmp[5634]*kernel[7]+tmp[5635]*kernel[8];
				ans[5535]<=tmp[5434]*kernel[0]+tmp[5435]*kernel[1]+tmp[5436]*kernel[2]+tmp[5534]*kernel[3]+tmp[5535]*kernel[4]+tmp[5536]*kernel[5]+tmp[5634]*kernel[6]+tmp[5635]*kernel[7]+tmp[5636]*kernel[8];
				ans[5536]<=tmp[5435]*kernel[0]+tmp[5436]*kernel[1]+tmp[5437]*kernel[2]+tmp[5535]*kernel[3]+tmp[5536]*kernel[4]+tmp[5537]*kernel[5]+tmp[5635]*kernel[6]+tmp[5636]*kernel[7]+tmp[5637]*kernel[8];
				ans[5537]<=tmp[5436]*kernel[0]+tmp[5437]*kernel[1]+tmp[5438]*kernel[2]+tmp[5536]*kernel[3]+tmp[5537]*kernel[4]+tmp[5538]*kernel[5]+tmp[5636]*kernel[6]+tmp[5637]*kernel[7]+tmp[5638]*kernel[8];
				ans[5538]<=tmp[5437]*kernel[0]+tmp[5438]*kernel[1]+tmp[5439]*kernel[2]+tmp[5537]*kernel[3]+tmp[5538]*kernel[4]+tmp[5539]*kernel[5]+tmp[5637]*kernel[6]+tmp[5638]*kernel[7]+tmp[5639]*kernel[8];
				ans[5539]<=tmp[5438]*kernel[0]+tmp[5439]*kernel[1]+tmp[5440]*kernel[2]+tmp[5538]*kernel[3]+tmp[5539]*kernel[4]+tmp[5540]*kernel[5]+tmp[5638]*kernel[6]+tmp[5639]*kernel[7]+tmp[5640]*kernel[8];
				ans[5540]<=tmp[5439]*kernel[0]+tmp[5440]*kernel[1]+tmp[5441]*kernel[2]+tmp[5539]*kernel[3]+tmp[5540]*kernel[4]+tmp[5541]*kernel[5]+tmp[5639]*kernel[6]+tmp[5640]*kernel[7]+tmp[5641]*kernel[8];
				ans[5541]<=tmp[5440]*kernel[0]+tmp[5441]*kernel[1]+tmp[5442]*kernel[2]+tmp[5540]*kernel[3]+tmp[5541]*kernel[4]+tmp[5542]*kernel[5]+tmp[5640]*kernel[6]+tmp[5641]*kernel[7]+tmp[5642]*kernel[8];
				ans[5542]<=tmp[5441]*kernel[0]+tmp[5442]*kernel[1]+tmp[5443]*kernel[2]+tmp[5541]*kernel[3]+tmp[5542]*kernel[4]+tmp[5543]*kernel[5]+tmp[5641]*kernel[6]+tmp[5642]*kernel[7]+tmp[5643]*kernel[8];
				ans[5543]<=tmp[5442]*kernel[0]+tmp[5443]*kernel[1]+tmp[5444]*kernel[2]+tmp[5542]*kernel[3]+tmp[5543]*kernel[4]+tmp[5544]*kernel[5]+tmp[5642]*kernel[6]+tmp[5643]*kernel[7]+tmp[5644]*kernel[8];
				ans[5544]<=tmp[5443]*kernel[0]+tmp[5444]*kernel[1]+tmp[5445]*kernel[2]+tmp[5543]*kernel[3]+tmp[5544]*kernel[4]+tmp[5545]*kernel[5]+tmp[5643]*kernel[6]+tmp[5644]*kernel[7]+tmp[5645]*kernel[8];
				ans[5545]<=tmp[5444]*kernel[0]+tmp[5445]*kernel[1]+tmp[5446]*kernel[2]+tmp[5544]*kernel[3]+tmp[5545]*kernel[4]+tmp[5546]*kernel[5]+tmp[5644]*kernel[6]+tmp[5645]*kernel[7]+tmp[5646]*kernel[8];
				ans[5546]<=tmp[5445]*kernel[0]+tmp[5446]*kernel[1]+tmp[5447]*kernel[2]+tmp[5545]*kernel[3]+tmp[5546]*kernel[4]+tmp[5547]*kernel[5]+tmp[5645]*kernel[6]+tmp[5646]*kernel[7]+tmp[5647]*kernel[8];
				ans[5547]<=tmp[5446]*kernel[0]+tmp[5447]*kernel[1]+tmp[5448]*kernel[2]+tmp[5546]*kernel[3]+tmp[5547]*kernel[4]+tmp[5548]*kernel[5]+tmp[5646]*kernel[6]+tmp[5647]*kernel[7]+tmp[5648]*kernel[8];
				ans[5548]<=tmp[5447]*kernel[0]+tmp[5448]*kernel[1]+tmp[5449]*kernel[2]+tmp[5547]*kernel[3]+tmp[5548]*kernel[4]+tmp[5549]*kernel[5]+tmp[5647]*kernel[6]+tmp[5648]*kernel[7]+tmp[5649]*kernel[8];
				ans[5549]<=tmp[5448]*kernel[0]+tmp[5449]*kernel[1]+tmp[5450]*kernel[2]+tmp[5548]*kernel[3]+tmp[5549]*kernel[4]+tmp[5550]*kernel[5]+tmp[5648]*kernel[6]+tmp[5649]*kernel[7]+tmp[5650]*kernel[8];
				ans[5550]<=tmp[5449]*kernel[0]+tmp[5450]*kernel[1]+tmp[5451]*kernel[2]+tmp[5549]*kernel[3]+tmp[5550]*kernel[4]+tmp[5551]*kernel[5]+tmp[5649]*kernel[6]+tmp[5650]*kernel[7]+tmp[5651]*kernel[8];
				ans[5551]<=tmp[5450]*kernel[0]+tmp[5451]*kernel[1]+tmp[5452]*kernel[2]+tmp[5550]*kernel[3]+tmp[5551]*kernel[4]+tmp[5552]*kernel[5]+tmp[5650]*kernel[6]+tmp[5651]*kernel[7]+tmp[5652]*kernel[8];
				ans[5552]<=tmp[5451]*kernel[0]+tmp[5452]*kernel[1]+tmp[5453]*kernel[2]+tmp[5551]*kernel[3]+tmp[5552]*kernel[4]+tmp[5553]*kernel[5]+tmp[5651]*kernel[6]+tmp[5652]*kernel[7]+tmp[5653]*kernel[8];
				ans[5553]<=tmp[5452]*kernel[0]+tmp[5453]*kernel[1]+tmp[5454]*kernel[2]+tmp[5552]*kernel[3]+tmp[5553]*kernel[4]+tmp[5554]*kernel[5]+tmp[5652]*kernel[6]+tmp[5653]*kernel[7]+tmp[5654]*kernel[8];
				ans[5554]<=tmp[5453]*kernel[0]+tmp[5454]*kernel[1]+tmp[5455]*kernel[2]+tmp[5553]*kernel[3]+tmp[5554]*kernel[4]+tmp[5555]*kernel[5]+tmp[5653]*kernel[6]+tmp[5654]*kernel[7]+tmp[5655]*kernel[8];
				ans[5555]<=tmp[5454]*kernel[0]+tmp[5455]*kernel[1]+tmp[5456]*kernel[2]+tmp[5554]*kernel[3]+tmp[5555]*kernel[4]+tmp[5556]*kernel[5]+tmp[5654]*kernel[6]+tmp[5655]*kernel[7]+tmp[5656]*kernel[8];
				ans[5556]<=tmp[5455]*kernel[0]+tmp[5456]*kernel[1]+tmp[5457]*kernel[2]+tmp[5555]*kernel[3]+tmp[5556]*kernel[4]+tmp[5557]*kernel[5]+tmp[5655]*kernel[6]+tmp[5656]*kernel[7]+tmp[5657]*kernel[8];
				ans[5557]<=tmp[5456]*kernel[0]+tmp[5457]*kernel[1]+tmp[5458]*kernel[2]+tmp[5556]*kernel[3]+tmp[5557]*kernel[4]+tmp[5558]*kernel[5]+tmp[5656]*kernel[6]+tmp[5657]*kernel[7]+tmp[5658]*kernel[8];
				ans[5558]<=tmp[5457]*kernel[0]+tmp[5458]*kernel[1]+tmp[5459]*kernel[2]+tmp[5557]*kernel[3]+tmp[5558]*kernel[4]+tmp[5559]*kernel[5]+tmp[5657]*kernel[6]+tmp[5658]*kernel[7]+tmp[5659]*kernel[8];
				ans[5559]<=tmp[5458]*kernel[0]+tmp[5459]*kernel[1]+tmp[5460]*kernel[2]+tmp[5558]*kernel[3]+tmp[5559]*kernel[4]+tmp[5560]*kernel[5]+tmp[5658]*kernel[6]+tmp[5659]*kernel[7]+tmp[5660]*kernel[8];
				ans[5560]<=tmp[5459]*kernel[0]+tmp[5460]*kernel[1]+tmp[5461]*kernel[2]+tmp[5559]*kernel[3]+tmp[5560]*kernel[4]+tmp[5561]*kernel[5]+tmp[5659]*kernel[6]+tmp[5660]*kernel[7]+tmp[5661]*kernel[8];
				ans[5561]<=tmp[5460]*kernel[0]+tmp[5461]*kernel[1]+tmp[5462]*kernel[2]+tmp[5560]*kernel[3]+tmp[5561]*kernel[4]+tmp[5562]*kernel[5]+tmp[5660]*kernel[6]+tmp[5661]*kernel[7]+tmp[5662]*kernel[8];
				ans[5562]<=tmp[5461]*kernel[0]+tmp[5462]*kernel[1]+tmp[5463]*kernel[2]+tmp[5561]*kernel[3]+tmp[5562]*kernel[4]+tmp[5563]*kernel[5]+tmp[5661]*kernel[6]+tmp[5662]*kernel[7]+tmp[5663]*kernel[8];
				ans[5563]<=tmp[5462]*kernel[0]+tmp[5463]*kernel[1]+tmp[5464]*kernel[2]+tmp[5562]*kernel[3]+tmp[5563]*kernel[4]+tmp[5564]*kernel[5]+tmp[5662]*kernel[6]+tmp[5663]*kernel[7]+tmp[5664]*kernel[8];
				ans[5564]<=tmp[5463]*kernel[0]+tmp[5464]*kernel[1]+tmp[5465]*kernel[2]+tmp[5563]*kernel[3]+tmp[5564]*kernel[4]+tmp[5565]*kernel[5]+tmp[5663]*kernel[6]+tmp[5664]*kernel[7]+tmp[5665]*kernel[8];
				ans[5565]<=tmp[5464]*kernel[0]+tmp[5465]*kernel[1]+tmp[5466]*kernel[2]+tmp[5564]*kernel[3]+tmp[5565]*kernel[4]+tmp[5566]*kernel[5]+tmp[5664]*kernel[6]+tmp[5665]*kernel[7]+tmp[5666]*kernel[8];
				ans[5566]<=tmp[5465]*kernel[0]+tmp[5466]*kernel[1]+tmp[5467]*kernel[2]+tmp[5565]*kernel[3]+tmp[5566]*kernel[4]+tmp[5567]*kernel[5]+tmp[5665]*kernel[6]+tmp[5666]*kernel[7]+tmp[5667]*kernel[8];
				ans[5567]<=tmp[5466]*kernel[0]+tmp[5467]*kernel[1]+tmp[5468]*kernel[2]+tmp[5566]*kernel[3]+tmp[5567]*kernel[4]+tmp[5568]*kernel[5]+tmp[5666]*kernel[6]+tmp[5667]*kernel[7]+tmp[5668]*kernel[8];
				ans[5568]<=tmp[5467]*kernel[0]+tmp[5468]*kernel[1]+tmp[5469]*kernel[2]+tmp[5567]*kernel[3]+tmp[5568]*kernel[4]+tmp[5569]*kernel[5]+tmp[5667]*kernel[6]+tmp[5668]*kernel[7]+tmp[5669]*kernel[8];
				ans[5569]<=tmp[5468]*kernel[0]+tmp[5469]*kernel[1]+tmp[5470]*kernel[2]+tmp[5568]*kernel[3]+tmp[5569]*kernel[4]+tmp[5570]*kernel[5]+tmp[5668]*kernel[6]+tmp[5669]*kernel[7]+tmp[5670]*kernel[8];
				ans[5570]<=tmp[5469]*kernel[0]+tmp[5470]*kernel[1]+tmp[5471]*kernel[2]+tmp[5569]*kernel[3]+tmp[5570]*kernel[4]+tmp[5571]*kernel[5]+tmp[5669]*kernel[6]+tmp[5670]*kernel[7]+tmp[5671]*kernel[8];
				ans[5571]<=tmp[5470]*kernel[0]+tmp[5471]*kernel[1]+tmp[5472]*kernel[2]+tmp[5570]*kernel[3]+tmp[5571]*kernel[4]+tmp[5572]*kernel[5]+tmp[5670]*kernel[6]+tmp[5671]*kernel[7]+tmp[5672]*kernel[8];
				ans[5572]<=tmp[5471]*kernel[0]+tmp[5472]*kernel[1]+tmp[5473]*kernel[2]+tmp[5571]*kernel[3]+tmp[5572]*kernel[4]+tmp[5573]*kernel[5]+tmp[5671]*kernel[6]+tmp[5672]*kernel[7]+tmp[5673]*kernel[8];
				ans[5573]<=tmp[5472]*kernel[0]+tmp[5473]*kernel[1]+tmp[5474]*kernel[2]+tmp[5572]*kernel[3]+tmp[5573]*kernel[4]+tmp[5574]*kernel[5]+tmp[5672]*kernel[6]+tmp[5673]*kernel[7]+tmp[5674]*kernel[8];
				ans[5574]<=tmp[5473]*kernel[0]+tmp[5474]*kernel[1]+tmp[5475]*kernel[2]+tmp[5573]*kernel[3]+tmp[5574]*kernel[4]+tmp[5575]*kernel[5]+tmp[5673]*kernel[6]+tmp[5674]*kernel[7]+tmp[5675]*kernel[8];
				ans[5575]<=tmp[5474]*kernel[0]+tmp[5475]*kernel[1]+tmp[5476]*kernel[2]+tmp[5574]*kernel[3]+tmp[5575]*kernel[4]+tmp[5576]*kernel[5]+tmp[5674]*kernel[6]+tmp[5675]*kernel[7]+tmp[5676]*kernel[8];
				ans[5576]<=tmp[5475]*kernel[0]+tmp[5476]*kernel[1]+tmp[5477]*kernel[2]+tmp[5575]*kernel[3]+tmp[5576]*kernel[4]+tmp[5577]*kernel[5]+tmp[5675]*kernel[6]+tmp[5676]*kernel[7]+tmp[5677]*kernel[8];
				ans[5577]<=tmp[5476]*kernel[0]+tmp[5477]*kernel[1]+tmp[5478]*kernel[2]+tmp[5576]*kernel[3]+tmp[5577]*kernel[4]+tmp[5578]*kernel[5]+tmp[5676]*kernel[6]+tmp[5677]*kernel[7]+tmp[5678]*kernel[8];
				ans[5578]<=tmp[5477]*kernel[0]+tmp[5478]*kernel[1]+tmp[5479]*kernel[2]+tmp[5577]*kernel[3]+tmp[5578]*kernel[4]+tmp[5579]*kernel[5]+tmp[5677]*kernel[6]+tmp[5678]*kernel[7]+tmp[5679]*kernel[8];
				ans[5579]<=tmp[5478]*kernel[0]+tmp[5479]*kernel[1]+tmp[5480]*kernel[2]+tmp[5578]*kernel[3]+tmp[5579]*kernel[4]+tmp[5580]*kernel[5]+tmp[5678]*kernel[6]+tmp[5679]*kernel[7]+tmp[5680]*kernel[8];
				ans[5580]<=tmp[5479]*kernel[0]+tmp[5480]*kernel[1]+tmp[5481]*kernel[2]+tmp[5579]*kernel[3]+tmp[5580]*kernel[4]+tmp[5581]*kernel[5]+tmp[5679]*kernel[6]+tmp[5680]*kernel[7]+tmp[5681]*kernel[8];
				ans[5581]<=tmp[5480]*kernel[0]+tmp[5481]*kernel[1]+tmp[5482]*kernel[2]+tmp[5580]*kernel[3]+tmp[5581]*kernel[4]+tmp[5582]*kernel[5]+tmp[5680]*kernel[6]+tmp[5681]*kernel[7]+tmp[5682]*kernel[8];
				ans[5582]<=tmp[5481]*kernel[0]+tmp[5482]*kernel[1]+tmp[5483]*kernel[2]+tmp[5581]*kernel[3]+tmp[5582]*kernel[4]+tmp[5583]*kernel[5]+tmp[5681]*kernel[6]+tmp[5682]*kernel[7]+tmp[5683]*kernel[8];
				ans[5583]<=tmp[5482]*kernel[0]+tmp[5483]*kernel[1]+tmp[5484]*kernel[2]+tmp[5582]*kernel[3]+tmp[5583]*kernel[4]+tmp[5584]*kernel[5]+tmp[5682]*kernel[6]+tmp[5683]*kernel[7]+tmp[5684]*kernel[8];
				ans[5584]<=tmp[5483]*kernel[0]+tmp[5484]*kernel[1]+tmp[5485]*kernel[2]+tmp[5583]*kernel[3]+tmp[5584]*kernel[4]+tmp[5585]*kernel[5]+tmp[5683]*kernel[6]+tmp[5684]*kernel[7]+tmp[5685]*kernel[8];
				ans[5585]<=tmp[5484]*kernel[0]+tmp[5485]*kernel[1]+tmp[5486]*kernel[2]+tmp[5584]*kernel[3]+tmp[5585]*kernel[4]+tmp[5586]*kernel[5]+tmp[5684]*kernel[6]+tmp[5685]*kernel[7]+tmp[5686]*kernel[8];
				ans[5586]<=tmp[5485]*kernel[0]+tmp[5486]*kernel[1]+tmp[5487]*kernel[2]+tmp[5585]*kernel[3]+tmp[5586]*kernel[4]+tmp[5587]*kernel[5]+tmp[5685]*kernel[6]+tmp[5686]*kernel[7]+tmp[5687]*kernel[8];
				ans[5587]<=tmp[5486]*kernel[0]+tmp[5487]*kernel[1]+tmp[5488]*kernel[2]+tmp[5586]*kernel[3]+tmp[5587]*kernel[4]+tmp[5588]*kernel[5]+tmp[5686]*kernel[6]+tmp[5687]*kernel[7]+tmp[5688]*kernel[8];
				ans[5588]<=tmp[5487]*kernel[0]+tmp[5488]*kernel[1]+tmp[5489]*kernel[2]+tmp[5587]*kernel[3]+tmp[5588]*kernel[4]+tmp[5589]*kernel[5]+tmp[5687]*kernel[6]+tmp[5688]*kernel[7]+tmp[5689]*kernel[8];
				ans[5589]<=tmp[5488]*kernel[0]+tmp[5489]*kernel[1]+tmp[5490]*kernel[2]+tmp[5588]*kernel[3]+tmp[5589]*kernel[4]+tmp[5590]*kernel[5]+tmp[5688]*kernel[6]+tmp[5689]*kernel[7]+tmp[5690]*kernel[8];
				ans[5590]<=tmp[5489]*kernel[0]+tmp[5490]*kernel[1]+tmp[5491]*kernel[2]+tmp[5589]*kernel[3]+tmp[5590]*kernel[4]+tmp[5591]*kernel[5]+tmp[5689]*kernel[6]+tmp[5690]*kernel[7]+tmp[5691]*kernel[8];
				ans[5591]<=tmp[5490]*kernel[0]+tmp[5491]*kernel[1]+tmp[5492]*kernel[2]+tmp[5590]*kernel[3]+tmp[5591]*kernel[4]+tmp[5592]*kernel[5]+tmp[5690]*kernel[6]+tmp[5691]*kernel[7]+tmp[5692]*kernel[8];
				ans[5592]<=tmp[5491]*kernel[0]+tmp[5492]*kernel[1]+tmp[5493]*kernel[2]+tmp[5591]*kernel[3]+tmp[5592]*kernel[4]+tmp[5593]*kernel[5]+tmp[5691]*kernel[6]+tmp[5692]*kernel[7]+tmp[5693]*kernel[8];
				ans[5593]<=tmp[5492]*kernel[0]+tmp[5493]*kernel[1]+tmp[5494]*kernel[2]+tmp[5592]*kernel[3]+tmp[5593]*kernel[4]+tmp[5594]*kernel[5]+tmp[5692]*kernel[6]+tmp[5693]*kernel[7]+tmp[5694]*kernel[8];
				ans[5594]<=tmp[5493]*kernel[0]+tmp[5494]*kernel[1]+tmp[5495]*kernel[2]+tmp[5593]*kernel[3]+tmp[5594]*kernel[4]+tmp[5595]*kernel[5]+tmp[5693]*kernel[6]+tmp[5694]*kernel[7]+tmp[5695]*kernel[8];
				ans[5595]<=tmp[5494]*kernel[0]+tmp[5495]*kernel[1]+tmp[5496]*kernel[2]+tmp[5594]*kernel[3]+tmp[5595]*kernel[4]+tmp[5596]*kernel[5]+tmp[5694]*kernel[6]+tmp[5695]*kernel[7]+tmp[5696]*kernel[8];
				ans[5596]<=tmp[5495]*kernel[0]+tmp[5496]*kernel[1]+tmp[5497]*kernel[2]+tmp[5595]*kernel[3]+tmp[5596]*kernel[4]+tmp[5597]*kernel[5]+tmp[5695]*kernel[6]+tmp[5696]*kernel[7]+tmp[5697]*kernel[8];
				ans[5597]<=tmp[5496]*kernel[0]+tmp[5497]*kernel[1]+tmp[5498]*kernel[2]+tmp[5596]*kernel[3]+tmp[5597]*kernel[4]+tmp[5598]*kernel[5]+tmp[5696]*kernel[6]+tmp[5697]*kernel[7]+tmp[5698]*kernel[8];
				ans[5598]<=tmp[5497]*kernel[0]+tmp[5498]*kernel[1]+tmp[5499]*kernel[2]+tmp[5597]*kernel[3]+tmp[5598]*kernel[4]+tmp[5599]*kernel[5]+tmp[5697]*kernel[6]+tmp[5698]*kernel[7]+tmp[5699]*kernel[8];
				ans[5599]<=tmp[5498]*kernel[0]+tmp[5499]*kernel[1]+tmp[5598]*kernel[3]+tmp[5599]*kernel[4]+tmp[5698]*kernel[6]+tmp[5699]*kernel[7];
				ans[5600]<=tmp[5500]*kernel[1]+tmp[5501]*kernel[2]+tmp[5600]*kernel[4]+tmp[5601]*kernel[5]+tmp[5700]*kernel[7]+tmp[5701]*kernel[8];
				ans[5601]<=tmp[5500]*kernel[0]+tmp[5501]*kernel[1]+tmp[5502]*kernel[2]+tmp[5600]*kernel[3]+tmp[5601]*kernel[4]+tmp[5602]*kernel[5]+tmp[5700]*kernel[6]+tmp[5701]*kernel[7]+tmp[5702]*kernel[8];
				ans[5602]<=tmp[5501]*kernel[0]+tmp[5502]*kernel[1]+tmp[5503]*kernel[2]+tmp[5601]*kernel[3]+tmp[5602]*kernel[4]+tmp[5603]*kernel[5]+tmp[5701]*kernel[6]+tmp[5702]*kernel[7]+tmp[5703]*kernel[8];
				ans[5603]<=tmp[5502]*kernel[0]+tmp[5503]*kernel[1]+tmp[5504]*kernel[2]+tmp[5602]*kernel[3]+tmp[5603]*kernel[4]+tmp[5604]*kernel[5]+tmp[5702]*kernel[6]+tmp[5703]*kernel[7]+tmp[5704]*kernel[8];
				ans[5604]<=tmp[5503]*kernel[0]+tmp[5504]*kernel[1]+tmp[5505]*kernel[2]+tmp[5603]*kernel[3]+tmp[5604]*kernel[4]+tmp[5605]*kernel[5]+tmp[5703]*kernel[6]+tmp[5704]*kernel[7]+tmp[5705]*kernel[8];
				ans[5605]<=tmp[5504]*kernel[0]+tmp[5505]*kernel[1]+tmp[5506]*kernel[2]+tmp[5604]*kernel[3]+tmp[5605]*kernel[4]+tmp[5606]*kernel[5]+tmp[5704]*kernel[6]+tmp[5705]*kernel[7]+tmp[5706]*kernel[8];
				ans[5606]<=tmp[5505]*kernel[0]+tmp[5506]*kernel[1]+tmp[5507]*kernel[2]+tmp[5605]*kernel[3]+tmp[5606]*kernel[4]+tmp[5607]*kernel[5]+tmp[5705]*kernel[6]+tmp[5706]*kernel[7]+tmp[5707]*kernel[8];
				ans[5607]<=tmp[5506]*kernel[0]+tmp[5507]*kernel[1]+tmp[5508]*kernel[2]+tmp[5606]*kernel[3]+tmp[5607]*kernel[4]+tmp[5608]*kernel[5]+tmp[5706]*kernel[6]+tmp[5707]*kernel[7]+tmp[5708]*kernel[8];
				ans[5608]<=tmp[5507]*kernel[0]+tmp[5508]*kernel[1]+tmp[5509]*kernel[2]+tmp[5607]*kernel[3]+tmp[5608]*kernel[4]+tmp[5609]*kernel[5]+tmp[5707]*kernel[6]+tmp[5708]*kernel[7]+tmp[5709]*kernel[8];
				ans[5609]<=tmp[5508]*kernel[0]+tmp[5509]*kernel[1]+tmp[5510]*kernel[2]+tmp[5608]*kernel[3]+tmp[5609]*kernel[4]+tmp[5610]*kernel[5]+tmp[5708]*kernel[6]+tmp[5709]*kernel[7]+tmp[5710]*kernel[8];
				ans[5610]<=tmp[5509]*kernel[0]+tmp[5510]*kernel[1]+tmp[5511]*kernel[2]+tmp[5609]*kernel[3]+tmp[5610]*kernel[4]+tmp[5611]*kernel[5]+tmp[5709]*kernel[6]+tmp[5710]*kernel[7]+tmp[5711]*kernel[8];
				ans[5611]<=tmp[5510]*kernel[0]+tmp[5511]*kernel[1]+tmp[5512]*kernel[2]+tmp[5610]*kernel[3]+tmp[5611]*kernel[4]+tmp[5612]*kernel[5]+tmp[5710]*kernel[6]+tmp[5711]*kernel[7]+tmp[5712]*kernel[8];
				ans[5612]<=tmp[5511]*kernel[0]+tmp[5512]*kernel[1]+tmp[5513]*kernel[2]+tmp[5611]*kernel[3]+tmp[5612]*kernel[4]+tmp[5613]*kernel[5]+tmp[5711]*kernel[6]+tmp[5712]*kernel[7]+tmp[5713]*kernel[8];
				ans[5613]<=tmp[5512]*kernel[0]+tmp[5513]*kernel[1]+tmp[5514]*kernel[2]+tmp[5612]*kernel[3]+tmp[5613]*kernel[4]+tmp[5614]*kernel[5]+tmp[5712]*kernel[6]+tmp[5713]*kernel[7]+tmp[5714]*kernel[8];
				ans[5614]<=tmp[5513]*kernel[0]+tmp[5514]*kernel[1]+tmp[5515]*kernel[2]+tmp[5613]*kernel[3]+tmp[5614]*kernel[4]+tmp[5615]*kernel[5]+tmp[5713]*kernel[6]+tmp[5714]*kernel[7]+tmp[5715]*kernel[8];
				ans[5615]<=tmp[5514]*kernel[0]+tmp[5515]*kernel[1]+tmp[5516]*kernel[2]+tmp[5614]*kernel[3]+tmp[5615]*kernel[4]+tmp[5616]*kernel[5]+tmp[5714]*kernel[6]+tmp[5715]*kernel[7]+tmp[5716]*kernel[8];
				ans[5616]<=tmp[5515]*kernel[0]+tmp[5516]*kernel[1]+tmp[5517]*kernel[2]+tmp[5615]*kernel[3]+tmp[5616]*kernel[4]+tmp[5617]*kernel[5]+tmp[5715]*kernel[6]+tmp[5716]*kernel[7]+tmp[5717]*kernel[8];
				ans[5617]<=tmp[5516]*kernel[0]+tmp[5517]*kernel[1]+tmp[5518]*kernel[2]+tmp[5616]*kernel[3]+tmp[5617]*kernel[4]+tmp[5618]*kernel[5]+tmp[5716]*kernel[6]+tmp[5717]*kernel[7]+tmp[5718]*kernel[8];
				ans[5618]<=tmp[5517]*kernel[0]+tmp[5518]*kernel[1]+tmp[5519]*kernel[2]+tmp[5617]*kernel[3]+tmp[5618]*kernel[4]+tmp[5619]*kernel[5]+tmp[5717]*kernel[6]+tmp[5718]*kernel[7]+tmp[5719]*kernel[8];
				ans[5619]<=tmp[5518]*kernel[0]+tmp[5519]*kernel[1]+tmp[5520]*kernel[2]+tmp[5618]*kernel[3]+tmp[5619]*kernel[4]+tmp[5620]*kernel[5]+tmp[5718]*kernel[6]+tmp[5719]*kernel[7]+tmp[5720]*kernel[8];
				ans[5620]<=tmp[5519]*kernel[0]+tmp[5520]*kernel[1]+tmp[5521]*kernel[2]+tmp[5619]*kernel[3]+tmp[5620]*kernel[4]+tmp[5621]*kernel[5]+tmp[5719]*kernel[6]+tmp[5720]*kernel[7]+tmp[5721]*kernel[8];
				ans[5621]<=tmp[5520]*kernel[0]+tmp[5521]*kernel[1]+tmp[5522]*kernel[2]+tmp[5620]*kernel[3]+tmp[5621]*kernel[4]+tmp[5622]*kernel[5]+tmp[5720]*kernel[6]+tmp[5721]*kernel[7]+tmp[5722]*kernel[8];
				ans[5622]<=tmp[5521]*kernel[0]+tmp[5522]*kernel[1]+tmp[5523]*kernel[2]+tmp[5621]*kernel[3]+tmp[5622]*kernel[4]+tmp[5623]*kernel[5]+tmp[5721]*kernel[6]+tmp[5722]*kernel[7]+tmp[5723]*kernel[8];
				ans[5623]<=tmp[5522]*kernel[0]+tmp[5523]*kernel[1]+tmp[5524]*kernel[2]+tmp[5622]*kernel[3]+tmp[5623]*kernel[4]+tmp[5624]*kernel[5]+tmp[5722]*kernel[6]+tmp[5723]*kernel[7]+tmp[5724]*kernel[8];
				ans[5624]<=tmp[5523]*kernel[0]+tmp[5524]*kernel[1]+tmp[5525]*kernel[2]+tmp[5623]*kernel[3]+tmp[5624]*kernel[4]+tmp[5625]*kernel[5]+tmp[5723]*kernel[6]+tmp[5724]*kernel[7]+tmp[5725]*kernel[8];
				ans[5625]<=tmp[5524]*kernel[0]+tmp[5525]*kernel[1]+tmp[5526]*kernel[2]+tmp[5624]*kernel[3]+tmp[5625]*kernel[4]+tmp[5626]*kernel[5]+tmp[5724]*kernel[6]+tmp[5725]*kernel[7]+tmp[5726]*kernel[8];
				ans[5626]<=tmp[5525]*kernel[0]+tmp[5526]*kernel[1]+tmp[5527]*kernel[2]+tmp[5625]*kernel[3]+tmp[5626]*kernel[4]+tmp[5627]*kernel[5]+tmp[5725]*kernel[6]+tmp[5726]*kernel[7]+tmp[5727]*kernel[8];
				ans[5627]<=tmp[5526]*kernel[0]+tmp[5527]*kernel[1]+tmp[5528]*kernel[2]+tmp[5626]*kernel[3]+tmp[5627]*kernel[4]+tmp[5628]*kernel[5]+tmp[5726]*kernel[6]+tmp[5727]*kernel[7]+tmp[5728]*kernel[8];
				ans[5628]<=tmp[5527]*kernel[0]+tmp[5528]*kernel[1]+tmp[5529]*kernel[2]+tmp[5627]*kernel[3]+tmp[5628]*kernel[4]+tmp[5629]*kernel[5]+tmp[5727]*kernel[6]+tmp[5728]*kernel[7]+tmp[5729]*kernel[8];
				ans[5629]<=tmp[5528]*kernel[0]+tmp[5529]*kernel[1]+tmp[5530]*kernel[2]+tmp[5628]*kernel[3]+tmp[5629]*kernel[4]+tmp[5630]*kernel[5]+tmp[5728]*kernel[6]+tmp[5729]*kernel[7]+tmp[5730]*kernel[8];
				ans[5630]<=tmp[5529]*kernel[0]+tmp[5530]*kernel[1]+tmp[5531]*kernel[2]+tmp[5629]*kernel[3]+tmp[5630]*kernel[4]+tmp[5631]*kernel[5]+tmp[5729]*kernel[6]+tmp[5730]*kernel[7]+tmp[5731]*kernel[8];
				ans[5631]<=tmp[5530]*kernel[0]+tmp[5531]*kernel[1]+tmp[5532]*kernel[2]+tmp[5630]*kernel[3]+tmp[5631]*kernel[4]+tmp[5632]*kernel[5]+tmp[5730]*kernel[6]+tmp[5731]*kernel[7]+tmp[5732]*kernel[8];
				ans[5632]<=tmp[5531]*kernel[0]+tmp[5532]*kernel[1]+tmp[5533]*kernel[2]+tmp[5631]*kernel[3]+tmp[5632]*kernel[4]+tmp[5633]*kernel[5]+tmp[5731]*kernel[6]+tmp[5732]*kernel[7]+tmp[5733]*kernel[8];
				ans[5633]<=tmp[5532]*kernel[0]+tmp[5533]*kernel[1]+tmp[5534]*kernel[2]+tmp[5632]*kernel[3]+tmp[5633]*kernel[4]+tmp[5634]*kernel[5]+tmp[5732]*kernel[6]+tmp[5733]*kernel[7]+tmp[5734]*kernel[8];
				ans[5634]<=tmp[5533]*kernel[0]+tmp[5534]*kernel[1]+tmp[5535]*kernel[2]+tmp[5633]*kernel[3]+tmp[5634]*kernel[4]+tmp[5635]*kernel[5]+tmp[5733]*kernel[6]+tmp[5734]*kernel[7]+tmp[5735]*kernel[8];
				ans[5635]<=tmp[5534]*kernel[0]+tmp[5535]*kernel[1]+tmp[5536]*kernel[2]+tmp[5634]*kernel[3]+tmp[5635]*kernel[4]+tmp[5636]*kernel[5]+tmp[5734]*kernel[6]+tmp[5735]*kernel[7]+tmp[5736]*kernel[8];
				ans[5636]<=tmp[5535]*kernel[0]+tmp[5536]*kernel[1]+tmp[5537]*kernel[2]+tmp[5635]*kernel[3]+tmp[5636]*kernel[4]+tmp[5637]*kernel[5]+tmp[5735]*kernel[6]+tmp[5736]*kernel[7]+tmp[5737]*kernel[8];
				ans[5637]<=tmp[5536]*kernel[0]+tmp[5537]*kernel[1]+tmp[5538]*kernel[2]+tmp[5636]*kernel[3]+tmp[5637]*kernel[4]+tmp[5638]*kernel[5]+tmp[5736]*kernel[6]+tmp[5737]*kernel[7]+tmp[5738]*kernel[8];
				ans[5638]<=tmp[5537]*kernel[0]+tmp[5538]*kernel[1]+tmp[5539]*kernel[2]+tmp[5637]*kernel[3]+tmp[5638]*kernel[4]+tmp[5639]*kernel[5]+tmp[5737]*kernel[6]+tmp[5738]*kernel[7]+tmp[5739]*kernel[8];
				ans[5639]<=tmp[5538]*kernel[0]+tmp[5539]*kernel[1]+tmp[5540]*kernel[2]+tmp[5638]*kernel[3]+tmp[5639]*kernel[4]+tmp[5640]*kernel[5]+tmp[5738]*kernel[6]+tmp[5739]*kernel[7]+tmp[5740]*kernel[8];
				ans[5640]<=tmp[5539]*kernel[0]+tmp[5540]*kernel[1]+tmp[5541]*kernel[2]+tmp[5639]*kernel[3]+tmp[5640]*kernel[4]+tmp[5641]*kernel[5]+tmp[5739]*kernel[6]+tmp[5740]*kernel[7]+tmp[5741]*kernel[8];
				ans[5641]<=tmp[5540]*kernel[0]+tmp[5541]*kernel[1]+tmp[5542]*kernel[2]+tmp[5640]*kernel[3]+tmp[5641]*kernel[4]+tmp[5642]*kernel[5]+tmp[5740]*kernel[6]+tmp[5741]*kernel[7]+tmp[5742]*kernel[8];
				ans[5642]<=tmp[5541]*kernel[0]+tmp[5542]*kernel[1]+tmp[5543]*kernel[2]+tmp[5641]*kernel[3]+tmp[5642]*kernel[4]+tmp[5643]*kernel[5]+tmp[5741]*kernel[6]+tmp[5742]*kernel[7]+tmp[5743]*kernel[8];
				ans[5643]<=tmp[5542]*kernel[0]+tmp[5543]*kernel[1]+tmp[5544]*kernel[2]+tmp[5642]*kernel[3]+tmp[5643]*kernel[4]+tmp[5644]*kernel[5]+tmp[5742]*kernel[6]+tmp[5743]*kernel[7]+tmp[5744]*kernel[8];
				ans[5644]<=tmp[5543]*kernel[0]+tmp[5544]*kernel[1]+tmp[5545]*kernel[2]+tmp[5643]*kernel[3]+tmp[5644]*kernel[4]+tmp[5645]*kernel[5]+tmp[5743]*kernel[6]+tmp[5744]*kernel[7]+tmp[5745]*kernel[8];
				ans[5645]<=tmp[5544]*kernel[0]+tmp[5545]*kernel[1]+tmp[5546]*kernel[2]+tmp[5644]*kernel[3]+tmp[5645]*kernel[4]+tmp[5646]*kernel[5]+tmp[5744]*kernel[6]+tmp[5745]*kernel[7]+tmp[5746]*kernel[8];
				ans[5646]<=tmp[5545]*kernel[0]+tmp[5546]*kernel[1]+tmp[5547]*kernel[2]+tmp[5645]*kernel[3]+tmp[5646]*kernel[4]+tmp[5647]*kernel[5]+tmp[5745]*kernel[6]+tmp[5746]*kernel[7]+tmp[5747]*kernel[8];
				ans[5647]<=tmp[5546]*kernel[0]+tmp[5547]*kernel[1]+tmp[5548]*kernel[2]+tmp[5646]*kernel[3]+tmp[5647]*kernel[4]+tmp[5648]*kernel[5]+tmp[5746]*kernel[6]+tmp[5747]*kernel[7]+tmp[5748]*kernel[8];
				ans[5648]<=tmp[5547]*kernel[0]+tmp[5548]*kernel[1]+tmp[5549]*kernel[2]+tmp[5647]*kernel[3]+tmp[5648]*kernel[4]+tmp[5649]*kernel[5]+tmp[5747]*kernel[6]+tmp[5748]*kernel[7]+tmp[5749]*kernel[8];
				ans[5649]<=tmp[5548]*kernel[0]+tmp[5549]*kernel[1]+tmp[5550]*kernel[2]+tmp[5648]*kernel[3]+tmp[5649]*kernel[4]+tmp[5650]*kernel[5]+tmp[5748]*kernel[6]+tmp[5749]*kernel[7]+tmp[5750]*kernel[8];
				ans[5650]<=tmp[5549]*kernel[0]+tmp[5550]*kernel[1]+tmp[5551]*kernel[2]+tmp[5649]*kernel[3]+tmp[5650]*kernel[4]+tmp[5651]*kernel[5]+tmp[5749]*kernel[6]+tmp[5750]*kernel[7]+tmp[5751]*kernel[8];
				ans[5651]<=tmp[5550]*kernel[0]+tmp[5551]*kernel[1]+tmp[5552]*kernel[2]+tmp[5650]*kernel[3]+tmp[5651]*kernel[4]+tmp[5652]*kernel[5]+tmp[5750]*kernel[6]+tmp[5751]*kernel[7]+tmp[5752]*kernel[8];
				ans[5652]<=tmp[5551]*kernel[0]+tmp[5552]*kernel[1]+tmp[5553]*kernel[2]+tmp[5651]*kernel[3]+tmp[5652]*kernel[4]+tmp[5653]*kernel[5]+tmp[5751]*kernel[6]+tmp[5752]*kernel[7]+tmp[5753]*kernel[8];
				ans[5653]<=tmp[5552]*kernel[0]+tmp[5553]*kernel[1]+tmp[5554]*kernel[2]+tmp[5652]*kernel[3]+tmp[5653]*kernel[4]+tmp[5654]*kernel[5]+tmp[5752]*kernel[6]+tmp[5753]*kernel[7]+tmp[5754]*kernel[8];
				ans[5654]<=tmp[5553]*kernel[0]+tmp[5554]*kernel[1]+tmp[5555]*kernel[2]+tmp[5653]*kernel[3]+tmp[5654]*kernel[4]+tmp[5655]*kernel[5]+tmp[5753]*kernel[6]+tmp[5754]*kernel[7]+tmp[5755]*kernel[8];
				ans[5655]<=tmp[5554]*kernel[0]+tmp[5555]*kernel[1]+tmp[5556]*kernel[2]+tmp[5654]*kernel[3]+tmp[5655]*kernel[4]+tmp[5656]*kernel[5]+tmp[5754]*kernel[6]+tmp[5755]*kernel[7]+tmp[5756]*kernel[8];
				ans[5656]<=tmp[5555]*kernel[0]+tmp[5556]*kernel[1]+tmp[5557]*kernel[2]+tmp[5655]*kernel[3]+tmp[5656]*kernel[4]+tmp[5657]*kernel[5]+tmp[5755]*kernel[6]+tmp[5756]*kernel[7]+tmp[5757]*kernel[8];
				ans[5657]<=tmp[5556]*kernel[0]+tmp[5557]*kernel[1]+tmp[5558]*kernel[2]+tmp[5656]*kernel[3]+tmp[5657]*kernel[4]+tmp[5658]*kernel[5]+tmp[5756]*kernel[6]+tmp[5757]*kernel[7]+tmp[5758]*kernel[8];
				ans[5658]<=tmp[5557]*kernel[0]+tmp[5558]*kernel[1]+tmp[5559]*kernel[2]+tmp[5657]*kernel[3]+tmp[5658]*kernel[4]+tmp[5659]*kernel[5]+tmp[5757]*kernel[6]+tmp[5758]*kernel[7]+tmp[5759]*kernel[8];
				ans[5659]<=tmp[5558]*kernel[0]+tmp[5559]*kernel[1]+tmp[5560]*kernel[2]+tmp[5658]*kernel[3]+tmp[5659]*kernel[4]+tmp[5660]*kernel[5]+tmp[5758]*kernel[6]+tmp[5759]*kernel[7]+tmp[5760]*kernel[8];
				ans[5660]<=tmp[5559]*kernel[0]+tmp[5560]*kernel[1]+tmp[5561]*kernel[2]+tmp[5659]*kernel[3]+tmp[5660]*kernel[4]+tmp[5661]*kernel[5]+tmp[5759]*kernel[6]+tmp[5760]*kernel[7]+tmp[5761]*kernel[8];
				ans[5661]<=tmp[5560]*kernel[0]+tmp[5561]*kernel[1]+tmp[5562]*kernel[2]+tmp[5660]*kernel[3]+tmp[5661]*kernel[4]+tmp[5662]*kernel[5]+tmp[5760]*kernel[6]+tmp[5761]*kernel[7]+tmp[5762]*kernel[8];
				ans[5662]<=tmp[5561]*kernel[0]+tmp[5562]*kernel[1]+tmp[5563]*kernel[2]+tmp[5661]*kernel[3]+tmp[5662]*kernel[4]+tmp[5663]*kernel[5]+tmp[5761]*kernel[6]+tmp[5762]*kernel[7]+tmp[5763]*kernel[8];
				ans[5663]<=tmp[5562]*kernel[0]+tmp[5563]*kernel[1]+tmp[5564]*kernel[2]+tmp[5662]*kernel[3]+tmp[5663]*kernel[4]+tmp[5664]*kernel[5]+tmp[5762]*kernel[6]+tmp[5763]*kernel[7]+tmp[5764]*kernel[8];
				ans[5664]<=tmp[5563]*kernel[0]+tmp[5564]*kernel[1]+tmp[5565]*kernel[2]+tmp[5663]*kernel[3]+tmp[5664]*kernel[4]+tmp[5665]*kernel[5]+tmp[5763]*kernel[6]+tmp[5764]*kernel[7]+tmp[5765]*kernel[8];
				ans[5665]<=tmp[5564]*kernel[0]+tmp[5565]*kernel[1]+tmp[5566]*kernel[2]+tmp[5664]*kernel[3]+tmp[5665]*kernel[4]+tmp[5666]*kernel[5]+tmp[5764]*kernel[6]+tmp[5765]*kernel[7]+tmp[5766]*kernel[8];
				ans[5666]<=tmp[5565]*kernel[0]+tmp[5566]*kernel[1]+tmp[5567]*kernel[2]+tmp[5665]*kernel[3]+tmp[5666]*kernel[4]+tmp[5667]*kernel[5]+tmp[5765]*kernel[6]+tmp[5766]*kernel[7]+tmp[5767]*kernel[8];
				ans[5667]<=tmp[5566]*kernel[0]+tmp[5567]*kernel[1]+tmp[5568]*kernel[2]+tmp[5666]*kernel[3]+tmp[5667]*kernel[4]+tmp[5668]*kernel[5]+tmp[5766]*kernel[6]+tmp[5767]*kernel[7]+tmp[5768]*kernel[8];
				ans[5668]<=tmp[5567]*kernel[0]+tmp[5568]*kernel[1]+tmp[5569]*kernel[2]+tmp[5667]*kernel[3]+tmp[5668]*kernel[4]+tmp[5669]*kernel[5]+tmp[5767]*kernel[6]+tmp[5768]*kernel[7]+tmp[5769]*kernel[8];
				ans[5669]<=tmp[5568]*kernel[0]+tmp[5569]*kernel[1]+tmp[5570]*kernel[2]+tmp[5668]*kernel[3]+tmp[5669]*kernel[4]+tmp[5670]*kernel[5]+tmp[5768]*kernel[6]+tmp[5769]*kernel[7]+tmp[5770]*kernel[8];
				ans[5670]<=tmp[5569]*kernel[0]+tmp[5570]*kernel[1]+tmp[5571]*kernel[2]+tmp[5669]*kernel[3]+tmp[5670]*kernel[4]+tmp[5671]*kernel[5]+tmp[5769]*kernel[6]+tmp[5770]*kernel[7]+tmp[5771]*kernel[8];
				ans[5671]<=tmp[5570]*kernel[0]+tmp[5571]*kernel[1]+tmp[5572]*kernel[2]+tmp[5670]*kernel[3]+tmp[5671]*kernel[4]+tmp[5672]*kernel[5]+tmp[5770]*kernel[6]+tmp[5771]*kernel[7]+tmp[5772]*kernel[8];
				ans[5672]<=tmp[5571]*kernel[0]+tmp[5572]*kernel[1]+tmp[5573]*kernel[2]+tmp[5671]*kernel[3]+tmp[5672]*kernel[4]+tmp[5673]*kernel[5]+tmp[5771]*kernel[6]+tmp[5772]*kernel[7]+tmp[5773]*kernel[8];
				ans[5673]<=tmp[5572]*kernel[0]+tmp[5573]*kernel[1]+tmp[5574]*kernel[2]+tmp[5672]*kernel[3]+tmp[5673]*kernel[4]+tmp[5674]*kernel[5]+tmp[5772]*kernel[6]+tmp[5773]*kernel[7]+tmp[5774]*kernel[8];
				ans[5674]<=tmp[5573]*kernel[0]+tmp[5574]*kernel[1]+tmp[5575]*kernel[2]+tmp[5673]*kernel[3]+tmp[5674]*kernel[4]+tmp[5675]*kernel[5]+tmp[5773]*kernel[6]+tmp[5774]*kernel[7]+tmp[5775]*kernel[8];
				ans[5675]<=tmp[5574]*kernel[0]+tmp[5575]*kernel[1]+tmp[5576]*kernel[2]+tmp[5674]*kernel[3]+tmp[5675]*kernel[4]+tmp[5676]*kernel[5]+tmp[5774]*kernel[6]+tmp[5775]*kernel[7]+tmp[5776]*kernel[8];
				ans[5676]<=tmp[5575]*kernel[0]+tmp[5576]*kernel[1]+tmp[5577]*kernel[2]+tmp[5675]*kernel[3]+tmp[5676]*kernel[4]+tmp[5677]*kernel[5]+tmp[5775]*kernel[6]+tmp[5776]*kernel[7]+tmp[5777]*kernel[8];
				ans[5677]<=tmp[5576]*kernel[0]+tmp[5577]*kernel[1]+tmp[5578]*kernel[2]+tmp[5676]*kernel[3]+tmp[5677]*kernel[4]+tmp[5678]*kernel[5]+tmp[5776]*kernel[6]+tmp[5777]*kernel[7]+tmp[5778]*kernel[8];
				ans[5678]<=tmp[5577]*kernel[0]+tmp[5578]*kernel[1]+tmp[5579]*kernel[2]+tmp[5677]*kernel[3]+tmp[5678]*kernel[4]+tmp[5679]*kernel[5]+tmp[5777]*kernel[6]+tmp[5778]*kernel[7]+tmp[5779]*kernel[8];
				ans[5679]<=tmp[5578]*kernel[0]+tmp[5579]*kernel[1]+tmp[5580]*kernel[2]+tmp[5678]*kernel[3]+tmp[5679]*kernel[4]+tmp[5680]*kernel[5]+tmp[5778]*kernel[6]+tmp[5779]*kernel[7]+tmp[5780]*kernel[8];
				ans[5680]<=tmp[5579]*kernel[0]+tmp[5580]*kernel[1]+tmp[5581]*kernel[2]+tmp[5679]*kernel[3]+tmp[5680]*kernel[4]+tmp[5681]*kernel[5]+tmp[5779]*kernel[6]+tmp[5780]*kernel[7]+tmp[5781]*kernel[8];
				ans[5681]<=tmp[5580]*kernel[0]+tmp[5581]*kernel[1]+tmp[5582]*kernel[2]+tmp[5680]*kernel[3]+tmp[5681]*kernel[4]+tmp[5682]*kernel[5]+tmp[5780]*kernel[6]+tmp[5781]*kernel[7]+tmp[5782]*kernel[8];
				ans[5682]<=tmp[5581]*kernel[0]+tmp[5582]*kernel[1]+tmp[5583]*kernel[2]+tmp[5681]*kernel[3]+tmp[5682]*kernel[4]+tmp[5683]*kernel[5]+tmp[5781]*kernel[6]+tmp[5782]*kernel[7]+tmp[5783]*kernel[8];
				ans[5683]<=tmp[5582]*kernel[0]+tmp[5583]*kernel[1]+tmp[5584]*kernel[2]+tmp[5682]*kernel[3]+tmp[5683]*kernel[4]+tmp[5684]*kernel[5]+tmp[5782]*kernel[6]+tmp[5783]*kernel[7]+tmp[5784]*kernel[8];
				ans[5684]<=tmp[5583]*kernel[0]+tmp[5584]*kernel[1]+tmp[5585]*kernel[2]+tmp[5683]*kernel[3]+tmp[5684]*kernel[4]+tmp[5685]*kernel[5]+tmp[5783]*kernel[6]+tmp[5784]*kernel[7]+tmp[5785]*kernel[8];
				ans[5685]<=tmp[5584]*kernel[0]+tmp[5585]*kernel[1]+tmp[5586]*kernel[2]+tmp[5684]*kernel[3]+tmp[5685]*kernel[4]+tmp[5686]*kernel[5]+tmp[5784]*kernel[6]+tmp[5785]*kernel[7]+tmp[5786]*kernel[8];
				ans[5686]<=tmp[5585]*kernel[0]+tmp[5586]*kernel[1]+tmp[5587]*kernel[2]+tmp[5685]*kernel[3]+tmp[5686]*kernel[4]+tmp[5687]*kernel[5]+tmp[5785]*kernel[6]+tmp[5786]*kernel[7]+tmp[5787]*kernel[8];
				ans[5687]<=tmp[5586]*kernel[0]+tmp[5587]*kernel[1]+tmp[5588]*kernel[2]+tmp[5686]*kernel[3]+tmp[5687]*kernel[4]+tmp[5688]*kernel[5]+tmp[5786]*kernel[6]+tmp[5787]*kernel[7]+tmp[5788]*kernel[8];
				ans[5688]<=tmp[5587]*kernel[0]+tmp[5588]*kernel[1]+tmp[5589]*kernel[2]+tmp[5687]*kernel[3]+tmp[5688]*kernel[4]+tmp[5689]*kernel[5]+tmp[5787]*kernel[6]+tmp[5788]*kernel[7]+tmp[5789]*kernel[8];
				ans[5689]<=tmp[5588]*kernel[0]+tmp[5589]*kernel[1]+tmp[5590]*kernel[2]+tmp[5688]*kernel[3]+tmp[5689]*kernel[4]+tmp[5690]*kernel[5]+tmp[5788]*kernel[6]+tmp[5789]*kernel[7]+tmp[5790]*kernel[8];
				ans[5690]<=tmp[5589]*kernel[0]+tmp[5590]*kernel[1]+tmp[5591]*kernel[2]+tmp[5689]*kernel[3]+tmp[5690]*kernel[4]+tmp[5691]*kernel[5]+tmp[5789]*kernel[6]+tmp[5790]*kernel[7]+tmp[5791]*kernel[8];
				ans[5691]<=tmp[5590]*kernel[0]+tmp[5591]*kernel[1]+tmp[5592]*kernel[2]+tmp[5690]*kernel[3]+tmp[5691]*kernel[4]+tmp[5692]*kernel[5]+tmp[5790]*kernel[6]+tmp[5791]*kernel[7]+tmp[5792]*kernel[8];
				ans[5692]<=tmp[5591]*kernel[0]+tmp[5592]*kernel[1]+tmp[5593]*kernel[2]+tmp[5691]*kernel[3]+tmp[5692]*kernel[4]+tmp[5693]*kernel[5]+tmp[5791]*kernel[6]+tmp[5792]*kernel[7]+tmp[5793]*kernel[8];
				ans[5693]<=tmp[5592]*kernel[0]+tmp[5593]*kernel[1]+tmp[5594]*kernel[2]+tmp[5692]*kernel[3]+tmp[5693]*kernel[4]+tmp[5694]*kernel[5]+tmp[5792]*kernel[6]+tmp[5793]*kernel[7]+tmp[5794]*kernel[8];
				ans[5694]<=tmp[5593]*kernel[0]+tmp[5594]*kernel[1]+tmp[5595]*kernel[2]+tmp[5693]*kernel[3]+tmp[5694]*kernel[4]+tmp[5695]*kernel[5]+tmp[5793]*kernel[6]+tmp[5794]*kernel[7]+tmp[5795]*kernel[8];
				ans[5695]<=tmp[5594]*kernel[0]+tmp[5595]*kernel[1]+tmp[5596]*kernel[2]+tmp[5694]*kernel[3]+tmp[5695]*kernel[4]+tmp[5696]*kernel[5]+tmp[5794]*kernel[6]+tmp[5795]*kernel[7]+tmp[5796]*kernel[8];
				ans[5696]<=tmp[5595]*kernel[0]+tmp[5596]*kernel[1]+tmp[5597]*kernel[2]+tmp[5695]*kernel[3]+tmp[5696]*kernel[4]+tmp[5697]*kernel[5]+tmp[5795]*kernel[6]+tmp[5796]*kernel[7]+tmp[5797]*kernel[8];
				ans[5697]<=tmp[5596]*kernel[0]+tmp[5597]*kernel[1]+tmp[5598]*kernel[2]+tmp[5696]*kernel[3]+tmp[5697]*kernel[4]+tmp[5698]*kernel[5]+tmp[5796]*kernel[6]+tmp[5797]*kernel[7]+tmp[5798]*kernel[8];
				ans[5698]<=tmp[5597]*kernel[0]+tmp[5598]*kernel[1]+tmp[5599]*kernel[2]+tmp[5697]*kernel[3]+tmp[5698]*kernel[4]+tmp[5699]*kernel[5]+tmp[5797]*kernel[6]+tmp[5798]*kernel[7]+tmp[5799]*kernel[8];
				ans[5699]<=tmp[5598]*kernel[0]+tmp[5599]*kernel[1]+tmp[5698]*kernel[3]+tmp[5699]*kernel[4]+tmp[5798]*kernel[6]+tmp[5799]*kernel[7];
				ans[5700]<=tmp[5600]*kernel[1]+tmp[5601]*kernel[2]+tmp[5700]*kernel[4]+tmp[5701]*kernel[5]+tmp[5800]*kernel[7]+tmp[5801]*kernel[8];
				ans[5701]<=tmp[5600]*kernel[0]+tmp[5601]*kernel[1]+tmp[5602]*kernel[2]+tmp[5700]*kernel[3]+tmp[5701]*kernel[4]+tmp[5702]*kernel[5]+tmp[5800]*kernel[6]+tmp[5801]*kernel[7]+tmp[5802]*kernel[8];
				ans[5702]<=tmp[5601]*kernel[0]+tmp[5602]*kernel[1]+tmp[5603]*kernel[2]+tmp[5701]*kernel[3]+tmp[5702]*kernel[4]+tmp[5703]*kernel[5]+tmp[5801]*kernel[6]+tmp[5802]*kernel[7]+tmp[5803]*kernel[8];
				ans[5703]<=tmp[5602]*kernel[0]+tmp[5603]*kernel[1]+tmp[5604]*kernel[2]+tmp[5702]*kernel[3]+tmp[5703]*kernel[4]+tmp[5704]*kernel[5]+tmp[5802]*kernel[6]+tmp[5803]*kernel[7]+tmp[5804]*kernel[8];
				ans[5704]<=tmp[5603]*kernel[0]+tmp[5604]*kernel[1]+tmp[5605]*kernel[2]+tmp[5703]*kernel[3]+tmp[5704]*kernel[4]+tmp[5705]*kernel[5]+tmp[5803]*kernel[6]+tmp[5804]*kernel[7]+tmp[5805]*kernel[8];
				ans[5705]<=tmp[5604]*kernel[0]+tmp[5605]*kernel[1]+tmp[5606]*kernel[2]+tmp[5704]*kernel[3]+tmp[5705]*kernel[4]+tmp[5706]*kernel[5]+tmp[5804]*kernel[6]+tmp[5805]*kernel[7]+tmp[5806]*kernel[8];
				ans[5706]<=tmp[5605]*kernel[0]+tmp[5606]*kernel[1]+tmp[5607]*kernel[2]+tmp[5705]*kernel[3]+tmp[5706]*kernel[4]+tmp[5707]*kernel[5]+tmp[5805]*kernel[6]+tmp[5806]*kernel[7]+tmp[5807]*kernel[8];
				ans[5707]<=tmp[5606]*kernel[0]+tmp[5607]*kernel[1]+tmp[5608]*kernel[2]+tmp[5706]*kernel[3]+tmp[5707]*kernel[4]+tmp[5708]*kernel[5]+tmp[5806]*kernel[6]+tmp[5807]*kernel[7]+tmp[5808]*kernel[8];
				ans[5708]<=tmp[5607]*kernel[0]+tmp[5608]*kernel[1]+tmp[5609]*kernel[2]+tmp[5707]*kernel[3]+tmp[5708]*kernel[4]+tmp[5709]*kernel[5]+tmp[5807]*kernel[6]+tmp[5808]*kernel[7]+tmp[5809]*kernel[8];
				ans[5709]<=tmp[5608]*kernel[0]+tmp[5609]*kernel[1]+tmp[5610]*kernel[2]+tmp[5708]*kernel[3]+tmp[5709]*kernel[4]+tmp[5710]*kernel[5]+tmp[5808]*kernel[6]+tmp[5809]*kernel[7]+tmp[5810]*kernel[8];
				ans[5710]<=tmp[5609]*kernel[0]+tmp[5610]*kernel[1]+tmp[5611]*kernel[2]+tmp[5709]*kernel[3]+tmp[5710]*kernel[4]+tmp[5711]*kernel[5]+tmp[5809]*kernel[6]+tmp[5810]*kernel[7]+tmp[5811]*kernel[8];
				ans[5711]<=tmp[5610]*kernel[0]+tmp[5611]*kernel[1]+tmp[5612]*kernel[2]+tmp[5710]*kernel[3]+tmp[5711]*kernel[4]+tmp[5712]*kernel[5]+tmp[5810]*kernel[6]+tmp[5811]*kernel[7]+tmp[5812]*kernel[8];
				ans[5712]<=tmp[5611]*kernel[0]+tmp[5612]*kernel[1]+tmp[5613]*kernel[2]+tmp[5711]*kernel[3]+tmp[5712]*kernel[4]+tmp[5713]*kernel[5]+tmp[5811]*kernel[6]+tmp[5812]*kernel[7]+tmp[5813]*kernel[8];
				ans[5713]<=tmp[5612]*kernel[0]+tmp[5613]*kernel[1]+tmp[5614]*kernel[2]+tmp[5712]*kernel[3]+tmp[5713]*kernel[4]+tmp[5714]*kernel[5]+tmp[5812]*kernel[6]+tmp[5813]*kernel[7]+tmp[5814]*kernel[8];
				ans[5714]<=tmp[5613]*kernel[0]+tmp[5614]*kernel[1]+tmp[5615]*kernel[2]+tmp[5713]*kernel[3]+tmp[5714]*kernel[4]+tmp[5715]*kernel[5]+tmp[5813]*kernel[6]+tmp[5814]*kernel[7]+tmp[5815]*kernel[8];
				ans[5715]<=tmp[5614]*kernel[0]+tmp[5615]*kernel[1]+tmp[5616]*kernel[2]+tmp[5714]*kernel[3]+tmp[5715]*kernel[4]+tmp[5716]*kernel[5]+tmp[5814]*kernel[6]+tmp[5815]*kernel[7]+tmp[5816]*kernel[8];
				ans[5716]<=tmp[5615]*kernel[0]+tmp[5616]*kernel[1]+tmp[5617]*kernel[2]+tmp[5715]*kernel[3]+tmp[5716]*kernel[4]+tmp[5717]*kernel[5]+tmp[5815]*kernel[6]+tmp[5816]*kernel[7]+tmp[5817]*kernel[8];
				ans[5717]<=tmp[5616]*kernel[0]+tmp[5617]*kernel[1]+tmp[5618]*kernel[2]+tmp[5716]*kernel[3]+tmp[5717]*kernel[4]+tmp[5718]*kernel[5]+tmp[5816]*kernel[6]+tmp[5817]*kernel[7]+tmp[5818]*kernel[8];
				ans[5718]<=tmp[5617]*kernel[0]+tmp[5618]*kernel[1]+tmp[5619]*kernel[2]+tmp[5717]*kernel[3]+tmp[5718]*kernel[4]+tmp[5719]*kernel[5]+tmp[5817]*kernel[6]+tmp[5818]*kernel[7]+tmp[5819]*kernel[8];
				ans[5719]<=tmp[5618]*kernel[0]+tmp[5619]*kernel[1]+tmp[5620]*kernel[2]+tmp[5718]*kernel[3]+tmp[5719]*kernel[4]+tmp[5720]*kernel[5]+tmp[5818]*kernel[6]+tmp[5819]*kernel[7]+tmp[5820]*kernel[8];
				ans[5720]<=tmp[5619]*kernel[0]+tmp[5620]*kernel[1]+tmp[5621]*kernel[2]+tmp[5719]*kernel[3]+tmp[5720]*kernel[4]+tmp[5721]*kernel[5]+tmp[5819]*kernel[6]+tmp[5820]*kernel[7]+tmp[5821]*kernel[8];
				ans[5721]<=tmp[5620]*kernel[0]+tmp[5621]*kernel[1]+tmp[5622]*kernel[2]+tmp[5720]*kernel[3]+tmp[5721]*kernel[4]+tmp[5722]*kernel[5]+tmp[5820]*kernel[6]+tmp[5821]*kernel[7]+tmp[5822]*kernel[8];
				ans[5722]<=tmp[5621]*kernel[0]+tmp[5622]*kernel[1]+tmp[5623]*kernel[2]+tmp[5721]*kernel[3]+tmp[5722]*kernel[4]+tmp[5723]*kernel[5]+tmp[5821]*kernel[6]+tmp[5822]*kernel[7]+tmp[5823]*kernel[8];
				ans[5723]<=tmp[5622]*kernel[0]+tmp[5623]*kernel[1]+tmp[5624]*kernel[2]+tmp[5722]*kernel[3]+tmp[5723]*kernel[4]+tmp[5724]*kernel[5]+tmp[5822]*kernel[6]+tmp[5823]*kernel[7]+tmp[5824]*kernel[8];
				ans[5724]<=tmp[5623]*kernel[0]+tmp[5624]*kernel[1]+tmp[5625]*kernel[2]+tmp[5723]*kernel[3]+tmp[5724]*kernel[4]+tmp[5725]*kernel[5]+tmp[5823]*kernel[6]+tmp[5824]*kernel[7]+tmp[5825]*kernel[8];
				ans[5725]<=tmp[5624]*kernel[0]+tmp[5625]*kernel[1]+tmp[5626]*kernel[2]+tmp[5724]*kernel[3]+tmp[5725]*kernel[4]+tmp[5726]*kernel[5]+tmp[5824]*kernel[6]+tmp[5825]*kernel[7]+tmp[5826]*kernel[8];
				ans[5726]<=tmp[5625]*kernel[0]+tmp[5626]*kernel[1]+tmp[5627]*kernel[2]+tmp[5725]*kernel[3]+tmp[5726]*kernel[4]+tmp[5727]*kernel[5]+tmp[5825]*kernel[6]+tmp[5826]*kernel[7]+tmp[5827]*kernel[8];
				ans[5727]<=tmp[5626]*kernel[0]+tmp[5627]*kernel[1]+tmp[5628]*kernel[2]+tmp[5726]*kernel[3]+tmp[5727]*kernel[4]+tmp[5728]*kernel[5]+tmp[5826]*kernel[6]+tmp[5827]*kernel[7]+tmp[5828]*kernel[8];
				ans[5728]<=tmp[5627]*kernel[0]+tmp[5628]*kernel[1]+tmp[5629]*kernel[2]+tmp[5727]*kernel[3]+tmp[5728]*kernel[4]+tmp[5729]*kernel[5]+tmp[5827]*kernel[6]+tmp[5828]*kernel[7]+tmp[5829]*kernel[8];
				ans[5729]<=tmp[5628]*kernel[0]+tmp[5629]*kernel[1]+tmp[5630]*kernel[2]+tmp[5728]*kernel[3]+tmp[5729]*kernel[4]+tmp[5730]*kernel[5]+tmp[5828]*kernel[6]+tmp[5829]*kernel[7]+tmp[5830]*kernel[8];
				ans[5730]<=tmp[5629]*kernel[0]+tmp[5630]*kernel[1]+tmp[5631]*kernel[2]+tmp[5729]*kernel[3]+tmp[5730]*kernel[4]+tmp[5731]*kernel[5]+tmp[5829]*kernel[6]+tmp[5830]*kernel[7]+tmp[5831]*kernel[8];
				ans[5731]<=tmp[5630]*kernel[0]+tmp[5631]*kernel[1]+tmp[5632]*kernel[2]+tmp[5730]*kernel[3]+tmp[5731]*kernel[4]+tmp[5732]*kernel[5]+tmp[5830]*kernel[6]+tmp[5831]*kernel[7]+tmp[5832]*kernel[8];
				ans[5732]<=tmp[5631]*kernel[0]+tmp[5632]*kernel[1]+tmp[5633]*kernel[2]+tmp[5731]*kernel[3]+tmp[5732]*kernel[4]+tmp[5733]*kernel[5]+tmp[5831]*kernel[6]+tmp[5832]*kernel[7]+tmp[5833]*kernel[8];
				ans[5733]<=tmp[5632]*kernel[0]+tmp[5633]*kernel[1]+tmp[5634]*kernel[2]+tmp[5732]*kernel[3]+tmp[5733]*kernel[4]+tmp[5734]*kernel[5]+tmp[5832]*kernel[6]+tmp[5833]*kernel[7]+tmp[5834]*kernel[8];
				ans[5734]<=tmp[5633]*kernel[0]+tmp[5634]*kernel[1]+tmp[5635]*kernel[2]+tmp[5733]*kernel[3]+tmp[5734]*kernel[4]+tmp[5735]*kernel[5]+tmp[5833]*kernel[6]+tmp[5834]*kernel[7]+tmp[5835]*kernel[8];
				ans[5735]<=tmp[5634]*kernel[0]+tmp[5635]*kernel[1]+tmp[5636]*kernel[2]+tmp[5734]*kernel[3]+tmp[5735]*kernel[4]+tmp[5736]*kernel[5]+tmp[5834]*kernel[6]+tmp[5835]*kernel[7]+tmp[5836]*kernel[8];
				ans[5736]<=tmp[5635]*kernel[0]+tmp[5636]*kernel[1]+tmp[5637]*kernel[2]+tmp[5735]*kernel[3]+tmp[5736]*kernel[4]+tmp[5737]*kernel[5]+tmp[5835]*kernel[6]+tmp[5836]*kernel[7]+tmp[5837]*kernel[8];
				ans[5737]<=tmp[5636]*kernel[0]+tmp[5637]*kernel[1]+tmp[5638]*kernel[2]+tmp[5736]*kernel[3]+tmp[5737]*kernel[4]+tmp[5738]*kernel[5]+tmp[5836]*kernel[6]+tmp[5837]*kernel[7]+tmp[5838]*kernel[8];
				ans[5738]<=tmp[5637]*kernel[0]+tmp[5638]*kernel[1]+tmp[5639]*kernel[2]+tmp[5737]*kernel[3]+tmp[5738]*kernel[4]+tmp[5739]*kernel[5]+tmp[5837]*kernel[6]+tmp[5838]*kernel[7]+tmp[5839]*kernel[8];
				ans[5739]<=tmp[5638]*kernel[0]+tmp[5639]*kernel[1]+tmp[5640]*kernel[2]+tmp[5738]*kernel[3]+tmp[5739]*kernel[4]+tmp[5740]*kernel[5]+tmp[5838]*kernel[6]+tmp[5839]*kernel[7]+tmp[5840]*kernel[8];
				ans[5740]<=tmp[5639]*kernel[0]+tmp[5640]*kernel[1]+tmp[5641]*kernel[2]+tmp[5739]*kernel[3]+tmp[5740]*kernel[4]+tmp[5741]*kernel[5]+tmp[5839]*kernel[6]+tmp[5840]*kernel[7]+tmp[5841]*kernel[8];
				ans[5741]<=tmp[5640]*kernel[0]+tmp[5641]*kernel[1]+tmp[5642]*kernel[2]+tmp[5740]*kernel[3]+tmp[5741]*kernel[4]+tmp[5742]*kernel[5]+tmp[5840]*kernel[6]+tmp[5841]*kernel[7]+tmp[5842]*kernel[8];
				ans[5742]<=tmp[5641]*kernel[0]+tmp[5642]*kernel[1]+tmp[5643]*kernel[2]+tmp[5741]*kernel[3]+tmp[5742]*kernel[4]+tmp[5743]*kernel[5]+tmp[5841]*kernel[6]+tmp[5842]*kernel[7]+tmp[5843]*kernel[8];
				ans[5743]<=tmp[5642]*kernel[0]+tmp[5643]*kernel[1]+tmp[5644]*kernel[2]+tmp[5742]*kernel[3]+tmp[5743]*kernel[4]+tmp[5744]*kernel[5]+tmp[5842]*kernel[6]+tmp[5843]*kernel[7]+tmp[5844]*kernel[8];
				ans[5744]<=tmp[5643]*kernel[0]+tmp[5644]*kernel[1]+tmp[5645]*kernel[2]+tmp[5743]*kernel[3]+tmp[5744]*kernel[4]+tmp[5745]*kernel[5]+tmp[5843]*kernel[6]+tmp[5844]*kernel[7]+tmp[5845]*kernel[8];
				ans[5745]<=tmp[5644]*kernel[0]+tmp[5645]*kernel[1]+tmp[5646]*kernel[2]+tmp[5744]*kernel[3]+tmp[5745]*kernel[4]+tmp[5746]*kernel[5]+tmp[5844]*kernel[6]+tmp[5845]*kernel[7]+tmp[5846]*kernel[8];
				ans[5746]<=tmp[5645]*kernel[0]+tmp[5646]*kernel[1]+tmp[5647]*kernel[2]+tmp[5745]*kernel[3]+tmp[5746]*kernel[4]+tmp[5747]*kernel[5]+tmp[5845]*kernel[6]+tmp[5846]*kernel[7]+tmp[5847]*kernel[8];
				ans[5747]<=tmp[5646]*kernel[0]+tmp[5647]*kernel[1]+tmp[5648]*kernel[2]+tmp[5746]*kernel[3]+tmp[5747]*kernel[4]+tmp[5748]*kernel[5]+tmp[5846]*kernel[6]+tmp[5847]*kernel[7]+tmp[5848]*kernel[8];
				ans[5748]<=tmp[5647]*kernel[0]+tmp[5648]*kernel[1]+tmp[5649]*kernel[2]+tmp[5747]*kernel[3]+tmp[5748]*kernel[4]+tmp[5749]*kernel[5]+tmp[5847]*kernel[6]+tmp[5848]*kernel[7]+tmp[5849]*kernel[8];
				ans[5749]<=tmp[5648]*kernel[0]+tmp[5649]*kernel[1]+tmp[5650]*kernel[2]+tmp[5748]*kernel[3]+tmp[5749]*kernel[4]+tmp[5750]*kernel[5]+tmp[5848]*kernel[6]+tmp[5849]*kernel[7]+tmp[5850]*kernel[8];
				ans[5750]<=tmp[5649]*kernel[0]+tmp[5650]*kernel[1]+tmp[5651]*kernel[2]+tmp[5749]*kernel[3]+tmp[5750]*kernel[4]+tmp[5751]*kernel[5]+tmp[5849]*kernel[6]+tmp[5850]*kernel[7]+tmp[5851]*kernel[8];
				ans[5751]<=tmp[5650]*kernel[0]+tmp[5651]*kernel[1]+tmp[5652]*kernel[2]+tmp[5750]*kernel[3]+tmp[5751]*kernel[4]+tmp[5752]*kernel[5]+tmp[5850]*kernel[6]+tmp[5851]*kernel[7]+tmp[5852]*kernel[8];
				ans[5752]<=tmp[5651]*kernel[0]+tmp[5652]*kernel[1]+tmp[5653]*kernel[2]+tmp[5751]*kernel[3]+tmp[5752]*kernel[4]+tmp[5753]*kernel[5]+tmp[5851]*kernel[6]+tmp[5852]*kernel[7]+tmp[5853]*kernel[8];
				ans[5753]<=tmp[5652]*kernel[0]+tmp[5653]*kernel[1]+tmp[5654]*kernel[2]+tmp[5752]*kernel[3]+tmp[5753]*kernel[4]+tmp[5754]*kernel[5]+tmp[5852]*kernel[6]+tmp[5853]*kernel[7]+tmp[5854]*kernel[8];
				ans[5754]<=tmp[5653]*kernel[0]+tmp[5654]*kernel[1]+tmp[5655]*kernel[2]+tmp[5753]*kernel[3]+tmp[5754]*kernel[4]+tmp[5755]*kernel[5]+tmp[5853]*kernel[6]+tmp[5854]*kernel[7]+tmp[5855]*kernel[8];
				ans[5755]<=tmp[5654]*kernel[0]+tmp[5655]*kernel[1]+tmp[5656]*kernel[2]+tmp[5754]*kernel[3]+tmp[5755]*kernel[4]+tmp[5756]*kernel[5]+tmp[5854]*kernel[6]+tmp[5855]*kernel[7]+tmp[5856]*kernel[8];
				ans[5756]<=tmp[5655]*kernel[0]+tmp[5656]*kernel[1]+tmp[5657]*kernel[2]+tmp[5755]*kernel[3]+tmp[5756]*kernel[4]+tmp[5757]*kernel[5]+tmp[5855]*kernel[6]+tmp[5856]*kernel[7]+tmp[5857]*kernel[8];
				ans[5757]<=tmp[5656]*kernel[0]+tmp[5657]*kernel[1]+tmp[5658]*kernel[2]+tmp[5756]*kernel[3]+tmp[5757]*kernel[4]+tmp[5758]*kernel[5]+tmp[5856]*kernel[6]+tmp[5857]*kernel[7]+tmp[5858]*kernel[8];
				ans[5758]<=tmp[5657]*kernel[0]+tmp[5658]*kernel[1]+tmp[5659]*kernel[2]+tmp[5757]*kernel[3]+tmp[5758]*kernel[4]+tmp[5759]*kernel[5]+tmp[5857]*kernel[6]+tmp[5858]*kernel[7]+tmp[5859]*kernel[8];
				ans[5759]<=tmp[5658]*kernel[0]+tmp[5659]*kernel[1]+tmp[5660]*kernel[2]+tmp[5758]*kernel[3]+tmp[5759]*kernel[4]+tmp[5760]*kernel[5]+tmp[5858]*kernel[6]+tmp[5859]*kernel[7]+tmp[5860]*kernel[8];
				ans[5760]<=tmp[5659]*kernel[0]+tmp[5660]*kernel[1]+tmp[5661]*kernel[2]+tmp[5759]*kernel[3]+tmp[5760]*kernel[4]+tmp[5761]*kernel[5]+tmp[5859]*kernel[6]+tmp[5860]*kernel[7]+tmp[5861]*kernel[8];
				ans[5761]<=tmp[5660]*kernel[0]+tmp[5661]*kernel[1]+tmp[5662]*kernel[2]+tmp[5760]*kernel[3]+tmp[5761]*kernel[4]+tmp[5762]*kernel[5]+tmp[5860]*kernel[6]+tmp[5861]*kernel[7]+tmp[5862]*kernel[8];
				ans[5762]<=tmp[5661]*kernel[0]+tmp[5662]*kernel[1]+tmp[5663]*kernel[2]+tmp[5761]*kernel[3]+tmp[5762]*kernel[4]+tmp[5763]*kernel[5]+tmp[5861]*kernel[6]+tmp[5862]*kernel[7]+tmp[5863]*kernel[8];
				ans[5763]<=tmp[5662]*kernel[0]+tmp[5663]*kernel[1]+tmp[5664]*kernel[2]+tmp[5762]*kernel[3]+tmp[5763]*kernel[4]+tmp[5764]*kernel[5]+tmp[5862]*kernel[6]+tmp[5863]*kernel[7]+tmp[5864]*kernel[8];
				ans[5764]<=tmp[5663]*kernel[0]+tmp[5664]*kernel[1]+tmp[5665]*kernel[2]+tmp[5763]*kernel[3]+tmp[5764]*kernel[4]+tmp[5765]*kernel[5]+tmp[5863]*kernel[6]+tmp[5864]*kernel[7]+tmp[5865]*kernel[8];
				ans[5765]<=tmp[5664]*kernel[0]+tmp[5665]*kernel[1]+tmp[5666]*kernel[2]+tmp[5764]*kernel[3]+tmp[5765]*kernel[4]+tmp[5766]*kernel[5]+tmp[5864]*kernel[6]+tmp[5865]*kernel[7]+tmp[5866]*kernel[8];
				ans[5766]<=tmp[5665]*kernel[0]+tmp[5666]*kernel[1]+tmp[5667]*kernel[2]+tmp[5765]*kernel[3]+tmp[5766]*kernel[4]+tmp[5767]*kernel[5]+tmp[5865]*kernel[6]+tmp[5866]*kernel[7]+tmp[5867]*kernel[8];
				ans[5767]<=tmp[5666]*kernel[0]+tmp[5667]*kernel[1]+tmp[5668]*kernel[2]+tmp[5766]*kernel[3]+tmp[5767]*kernel[4]+tmp[5768]*kernel[5]+tmp[5866]*kernel[6]+tmp[5867]*kernel[7]+tmp[5868]*kernel[8];
				ans[5768]<=tmp[5667]*kernel[0]+tmp[5668]*kernel[1]+tmp[5669]*kernel[2]+tmp[5767]*kernel[3]+tmp[5768]*kernel[4]+tmp[5769]*kernel[5]+tmp[5867]*kernel[6]+tmp[5868]*kernel[7]+tmp[5869]*kernel[8];
				ans[5769]<=tmp[5668]*kernel[0]+tmp[5669]*kernel[1]+tmp[5670]*kernel[2]+tmp[5768]*kernel[3]+tmp[5769]*kernel[4]+tmp[5770]*kernel[5]+tmp[5868]*kernel[6]+tmp[5869]*kernel[7]+tmp[5870]*kernel[8];
				ans[5770]<=tmp[5669]*kernel[0]+tmp[5670]*kernel[1]+tmp[5671]*kernel[2]+tmp[5769]*kernel[3]+tmp[5770]*kernel[4]+tmp[5771]*kernel[5]+tmp[5869]*kernel[6]+tmp[5870]*kernel[7]+tmp[5871]*kernel[8];
				ans[5771]<=tmp[5670]*kernel[0]+tmp[5671]*kernel[1]+tmp[5672]*kernel[2]+tmp[5770]*kernel[3]+tmp[5771]*kernel[4]+tmp[5772]*kernel[5]+tmp[5870]*kernel[6]+tmp[5871]*kernel[7]+tmp[5872]*kernel[8];
				ans[5772]<=tmp[5671]*kernel[0]+tmp[5672]*kernel[1]+tmp[5673]*kernel[2]+tmp[5771]*kernel[3]+tmp[5772]*kernel[4]+tmp[5773]*kernel[5]+tmp[5871]*kernel[6]+tmp[5872]*kernel[7]+tmp[5873]*kernel[8];
				ans[5773]<=tmp[5672]*kernel[0]+tmp[5673]*kernel[1]+tmp[5674]*kernel[2]+tmp[5772]*kernel[3]+tmp[5773]*kernel[4]+tmp[5774]*kernel[5]+tmp[5872]*kernel[6]+tmp[5873]*kernel[7]+tmp[5874]*kernel[8];
				ans[5774]<=tmp[5673]*kernel[0]+tmp[5674]*kernel[1]+tmp[5675]*kernel[2]+tmp[5773]*kernel[3]+tmp[5774]*kernel[4]+tmp[5775]*kernel[5]+tmp[5873]*kernel[6]+tmp[5874]*kernel[7]+tmp[5875]*kernel[8];
				ans[5775]<=tmp[5674]*kernel[0]+tmp[5675]*kernel[1]+tmp[5676]*kernel[2]+tmp[5774]*kernel[3]+tmp[5775]*kernel[4]+tmp[5776]*kernel[5]+tmp[5874]*kernel[6]+tmp[5875]*kernel[7]+tmp[5876]*kernel[8];
				ans[5776]<=tmp[5675]*kernel[0]+tmp[5676]*kernel[1]+tmp[5677]*kernel[2]+tmp[5775]*kernel[3]+tmp[5776]*kernel[4]+tmp[5777]*kernel[5]+tmp[5875]*kernel[6]+tmp[5876]*kernel[7]+tmp[5877]*kernel[8];
				ans[5777]<=tmp[5676]*kernel[0]+tmp[5677]*kernel[1]+tmp[5678]*kernel[2]+tmp[5776]*kernel[3]+tmp[5777]*kernel[4]+tmp[5778]*kernel[5]+tmp[5876]*kernel[6]+tmp[5877]*kernel[7]+tmp[5878]*kernel[8];
				ans[5778]<=tmp[5677]*kernel[0]+tmp[5678]*kernel[1]+tmp[5679]*kernel[2]+tmp[5777]*kernel[3]+tmp[5778]*kernel[4]+tmp[5779]*kernel[5]+tmp[5877]*kernel[6]+tmp[5878]*kernel[7]+tmp[5879]*kernel[8];
				ans[5779]<=tmp[5678]*kernel[0]+tmp[5679]*kernel[1]+tmp[5680]*kernel[2]+tmp[5778]*kernel[3]+tmp[5779]*kernel[4]+tmp[5780]*kernel[5]+tmp[5878]*kernel[6]+tmp[5879]*kernel[7]+tmp[5880]*kernel[8];
				ans[5780]<=tmp[5679]*kernel[0]+tmp[5680]*kernel[1]+tmp[5681]*kernel[2]+tmp[5779]*kernel[3]+tmp[5780]*kernel[4]+tmp[5781]*kernel[5]+tmp[5879]*kernel[6]+tmp[5880]*kernel[7]+tmp[5881]*kernel[8];
				ans[5781]<=tmp[5680]*kernel[0]+tmp[5681]*kernel[1]+tmp[5682]*kernel[2]+tmp[5780]*kernel[3]+tmp[5781]*kernel[4]+tmp[5782]*kernel[5]+tmp[5880]*kernel[6]+tmp[5881]*kernel[7]+tmp[5882]*kernel[8];
				ans[5782]<=tmp[5681]*kernel[0]+tmp[5682]*kernel[1]+tmp[5683]*kernel[2]+tmp[5781]*kernel[3]+tmp[5782]*kernel[4]+tmp[5783]*kernel[5]+tmp[5881]*kernel[6]+tmp[5882]*kernel[7]+tmp[5883]*kernel[8];
				ans[5783]<=tmp[5682]*kernel[0]+tmp[5683]*kernel[1]+tmp[5684]*kernel[2]+tmp[5782]*kernel[3]+tmp[5783]*kernel[4]+tmp[5784]*kernel[5]+tmp[5882]*kernel[6]+tmp[5883]*kernel[7]+tmp[5884]*kernel[8];
				ans[5784]<=tmp[5683]*kernel[0]+tmp[5684]*kernel[1]+tmp[5685]*kernel[2]+tmp[5783]*kernel[3]+tmp[5784]*kernel[4]+tmp[5785]*kernel[5]+tmp[5883]*kernel[6]+tmp[5884]*kernel[7]+tmp[5885]*kernel[8];
				ans[5785]<=tmp[5684]*kernel[0]+tmp[5685]*kernel[1]+tmp[5686]*kernel[2]+tmp[5784]*kernel[3]+tmp[5785]*kernel[4]+tmp[5786]*kernel[5]+tmp[5884]*kernel[6]+tmp[5885]*kernel[7]+tmp[5886]*kernel[8];
				ans[5786]<=tmp[5685]*kernel[0]+tmp[5686]*kernel[1]+tmp[5687]*kernel[2]+tmp[5785]*kernel[3]+tmp[5786]*kernel[4]+tmp[5787]*kernel[5]+tmp[5885]*kernel[6]+tmp[5886]*kernel[7]+tmp[5887]*kernel[8];
				ans[5787]<=tmp[5686]*kernel[0]+tmp[5687]*kernel[1]+tmp[5688]*kernel[2]+tmp[5786]*kernel[3]+tmp[5787]*kernel[4]+tmp[5788]*kernel[5]+tmp[5886]*kernel[6]+tmp[5887]*kernel[7]+tmp[5888]*kernel[8];
				ans[5788]<=tmp[5687]*kernel[0]+tmp[5688]*kernel[1]+tmp[5689]*kernel[2]+tmp[5787]*kernel[3]+tmp[5788]*kernel[4]+tmp[5789]*kernel[5]+tmp[5887]*kernel[6]+tmp[5888]*kernel[7]+tmp[5889]*kernel[8];
				ans[5789]<=tmp[5688]*kernel[0]+tmp[5689]*kernel[1]+tmp[5690]*kernel[2]+tmp[5788]*kernel[3]+tmp[5789]*kernel[4]+tmp[5790]*kernel[5]+tmp[5888]*kernel[6]+tmp[5889]*kernel[7]+tmp[5890]*kernel[8];
				ans[5790]<=tmp[5689]*kernel[0]+tmp[5690]*kernel[1]+tmp[5691]*kernel[2]+tmp[5789]*kernel[3]+tmp[5790]*kernel[4]+tmp[5791]*kernel[5]+tmp[5889]*kernel[6]+tmp[5890]*kernel[7]+tmp[5891]*kernel[8];
				ans[5791]<=tmp[5690]*kernel[0]+tmp[5691]*kernel[1]+tmp[5692]*kernel[2]+tmp[5790]*kernel[3]+tmp[5791]*kernel[4]+tmp[5792]*kernel[5]+tmp[5890]*kernel[6]+tmp[5891]*kernel[7]+tmp[5892]*kernel[8];
				ans[5792]<=tmp[5691]*kernel[0]+tmp[5692]*kernel[1]+tmp[5693]*kernel[2]+tmp[5791]*kernel[3]+tmp[5792]*kernel[4]+tmp[5793]*kernel[5]+tmp[5891]*kernel[6]+tmp[5892]*kernel[7]+tmp[5893]*kernel[8];
				ans[5793]<=tmp[5692]*kernel[0]+tmp[5693]*kernel[1]+tmp[5694]*kernel[2]+tmp[5792]*kernel[3]+tmp[5793]*kernel[4]+tmp[5794]*kernel[5]+tmp[5892]*kernel[6]+tmp[5893]*kernel[7]+tmp[5894]*kernel[8];
				ans[5794]<=tmp[5693]*kernel[0]+tmp[5694]*kernel[1]+tmp[5695]*kernel[2]+tmp[5793]*kernel[3]+tmp[5794]*kernel[4]+tmp[5795]*kernel[5]+tmp[5893]*kernel[6]+tmp[5894]*kernel[7]+tmp[5895]*kernel[8];
				ans[5795]<=tmp[5694]*kernel[0]+tmp[5695]*kernel[1]+tmp[5696]*kernel[2]+tmp[5794]*kernel[3]+tmp[5795]*kernel[4]+tmp[5796]*kernel[5]+tmp[5894]*kernel[6]+tmp[5895]*kernel[7]+tmp[5896]*kernel[8];
				ans[5796]<=tmp[5695]*kernel[0]+tmp[5696]*kernel[1]+tmp[5697]*kernel[2]+tmp[5795]*kernel[3]+tmp[5796]*kernel[4]+tmp[5797]*kernel[5]+tmp[5895]*kernel[6]+tmp[5896]*kernel[7]+tmp[5897]*kernel[8];
				ans[5797]<=tmp[5696]*kernel[0]+tmp[5697]*kernel[1]+tmp[5698]*kernel[2]+tmp[5796]*kernel[3]+tmp[5797]*kernel[4]+tmp[5798]*kernel[5]+tmp[5896]*kernel[6]+tmp[5897]*kernel[7]+tmp[5898]*kernel[8];
				ans[5798]<=tmp[5697]*kernel[0]+tmp[5698]*kernel[1]+tmp[5699]*kernel[2]+tmp[5797]*kernel[3]+tmp[5798]*kernel[4]+tmp[5799]*kernel[5]+tmp[5897]*kernel[6]+tmp[5898]*kernel[7]+tmp[5899]*kernel[8];
				ans[5799]<=tmp[5698]*kernel[0]+tmp[5699]*kernel[1]+tmp[5798]*kernel[3]+tmp[5799]*kernel[4]+tmp[5898]*kernel[6]+tmp[5899]*kernel[7];
				ans[5800]<=tmp[5700]*kernel[1]+tmp[5701]*kernel[2]+tmp[5800]*kernel[4]+tmp[5801]*kernel[5]+tmp[5900]*kernel[7]+tmp[5901]*kernel[8];
				ans[5801]<=tmp[5700]*kernel[0]+tmp[5701]*kernel[1]+tmp[5702]*kernel[2]+tmp[5800]*kernel[3]+tmp[5801]*kernel[4]+tmp[5802]*kernel[5]+tmp[5900]*kernel[6]+tmp[5901]*kernel[7]+tmp[5902]*kernel[8];
				ans[5802]<=tmp[5701]*kernel[0]+tmp[5702]*kernel[1]+tmp[5703]*kernel[2]+tmp[5801]*kernel[3]+tmp[5802]*kernel[4]+tmp[5803]*kernel[5]+tmp[5901]*kernel[6]+tmp[5902]*kernel[7]+tmp[5903]*kernel[8];
				ans[5803]<=tmp[5702]*kernel[0]+tmp[5703]*kernel[1]+tmp[5704]*kernel[2]+tmp[5802]*kernel[3]+tmp[5803]*kernel[4]+tmp[5804]*kernel[5]+tmp[5902]*kernel[6]+tmp[5903]*kernel[7]+tmp[5904]*kernel[8];
				ans[5804]<=tmp[5703]*kernel[0]+tmp[5704]*kernel[1]+tmp[5705]*kernel[2]+tmp[5803]*kernel[3]+tmp[5804]*kernel[4]+tmp[5805]*kernel[5]+tmp[5903]*kernel[6]+tmp[5904]*kernel[7]+tmp[5905]*kernel[8];
				ans[5805]<=tmp[5704]*kernel[0]+tmp[5705]*kernel[1]+tmp[5706]*kernel[2]+tmp[5804]*kernel[3]+tmp[5805]*kernel[4]+tmp[5806]*kernel[5]+tmp[5904]*kernel[6]+tmp[5905]*kernel[7]+tmp[5906]*kernel[8];
				ans[5806]<=tmp[5705]*kernel[0]+tmp[5706]*kernel[1]+tmp[5707]*kernel[2]+tmp[5805]*kernel[3]+tmp[5806]*kernel[4]+tmp[5807]*kernel[5]+tmp[5905]*kernel[6]+tmp[5906]*kernel[7]+tmp[5907]*kernel[8];
				ans[5807]<=tmp[5706]*kernel[0]+tmp[5707]*kernel[1]+tmp[5708]*kernel[2]+tmp[5806]*kernel[3]+tmp[5807]*kernel[4]+tmp[5808]*kernel[5]+tmp[5906]*kernel[6]+tmp[5907]*kernel[7]+tmp[5908]*kernel[8];
				ans[5808]<=tmp[5707]*kernel[0]+tmp[5708]*kernel[1]+tmp[5709]*kernel[2]+tmp[5807]*kernel[3]+tmp[5808]*kernel[4]+tmp[5809]*kernel[5]+tmp[5907]*kernel[6]+tmp[5908]*kernel[7]+tmp[5909]*kernel[8];
				ans[5809]<=tmp[5708]*kernel[0]+tmp[5709]*kernel[1]+tmp[5710]*kernel[2]+tmp[5808]*kernel[3]+tmp[5809]*kernel[4]+tmp[5810]*kernel[5]+tmp[5908]*kernel[6]+tmp[5909]*kernel[7]+tmp[5910]*kernel[8];
				ans[5810]<=tmp[5709]*kernel[0]+tmp[5710]*kernel[1]+tmp[5711]*kernel[2]+tmp[5809]*kernel[3]+tmp[5810]*kernel[4]+tmp[5811]*kernel[5]+tmp[5909]*kernel[6]+tmp[5910]*kernel[7]+tmp[5911]*kernel[8];
				ans[5811]<=tmp[5710]*kernel[0]+tmp[5711]*kernel[1]+tmp[5712]*kernel[2]+tmp[5810]*kernel[3]+tmp[5811]*kernel[4]+tmp[5812]*kernel[5]+tmp[5910]*kernel[6]+tmp[5911]*kernel[7]+tmp[5912]*kernel[8];
				ans[5812]<=tmp[5711]*kernel[0]+tmp[5712]*kernel[1]+tmp[5713]*kernel[2]+tmp[5811]*kernel[3]+tmp[5812]*kernel[4]+tmp[5813]*kernel[5]+tmp[5911]*kernel[6]+tmp[5912]*kernel[7]+tmp[5913]*kernel[8];
				ans[5813]<=tmp[5712]*kernel[0]+tmp[5713]*kernel[1]+tmp[5714]*kernel[2]+tmp[5812]*kernel[3]+tmp[5813]*kernel[4]+tmp[5814]*kernel[5]+tmp[5912]*kernel[6]+tmp[5913]*kernel[7]+tmp[5914]*kernel[8];
				ans[5814]<=tmp[5713]*kernel[0]+tmp[5714]*kernel[1]+tmp[5715]*kernel[2]+tmp[5813]*kernel[3]+tmp[5814]*kernel[4]+tmp[5815]*kernel[5]+tmp[5913]*kernel[6]+tmp[5914]*kernel[7]+tmp[5915]*kernel[8];
				ans[5815]<=tmp[5714]*kernel[0]+tmp[5715]*kernel[1]+tmp[5716]*kernel[2]+tmp[5814]*kernel[3]+tmp[5815]*kernel[4]+tmp[5816]*kernel[5]+tmp[5914]*kernel[6]+tmp[5915]*kernel[7]+tmp[5916]*kernel[8];
				ans[5816]<=tmp[5715]*kernel[0]+tmp[5716]*kernel[1]+tmp[5717]*kernel[2]+tmp[5815]*kernel[3]+tmp[5816]*kernel[4]+tmp[5817]*kernel[5]+tmp[5915]*kernel[6]+tmp[5916]*kernel[7]+tmp[5917]*kernel[8];
				ans[5817]<=tmp[5716]*kernel[0]+tmp[5717]*kernel[1]+tmp[5718]*kernel[2]+tmp[5816]*kernel[3]+tmp[5817]*kernel[4]+tmp[5818]*kernel[5]+tmp[5916]*kernel[6]+tmp[5917]*kernel[7]+tmp[5918]*kernel[8];
				ans[5818]<=tmp[5717]*kernel[0]+tmp[5718]*kernel[1]+tmp[5719]*kernel[2]+tmp[5817]*kernel[3]+tmp[5818]*kernel[4]+tmp[5819]*kernel[5]+tmp[5917]*kernel[6]+tmp[5918]*kernel[7]+tmp[5919]*kernel[8];
				ans[5819]<=tmp[5718]*kernel[0]+tmp[5719]*kernel[1]+tmp[5720]*kernel[2]+tmp[5818]*kernel[3]+tmp[5819]*kernel[4]+tmp[5820]*kernel[5]+tmp[5918]*kernel[6]+tmp[5919]*kernel[7]+tmp[5920]*kernel[8];
				ans[5820]<=tmp[5719]*kernel[0]+tmp[5720]*kernel[1]+tmp[5721]*kernel[2]+tmp[5819]*kernel[3]+tmp[5820]*kernel[4]+tmp[5821]*kernel[5]+tmp[5919]*kernel[6]+tmp[5920]*kernel[7]+tmp[5921]*kernel[8];
				ans[5821]<=tmp[5720]*kernel[0]+tmp[5721]*kernel[1]+tmp[5722]*kernel[2]+tmp[5820]*kernel[3]+tmp[5821]*kernel[4]+tmp[5822]*kernel[5]+tmp[5920]*kernel[6]+tmp[5921]*kernel[7]+tmp[5922]*kernel[8];
				ans[5822]<=tmp[5721]*kernel[0]+tmp[5722]*kernel[1]+tmp[5723]*kernel[2]+tmp[5821]*kernel[3]+tmp[5822]*kernel[4]+tmp[5823]*kernel[5]+tmp[5921]*kernel[6]+tmp[5922]*kernel[7]+tmp[5923]*kernel[8];
				ans[5823]<=tmp[5722]*kernel[0]+tmp[5723]*kernel[1]+tmp[5724]*kernel[2]+tmp[5822]*kernel[3]+tmp[5823]*kernel[4]+tmp[5824]*kernel[5]+tmp[5922]*kernel[6]+tmp[5923]*kernel[7]+tmp[5924]*kernel[8];
				ans[5824]<=tmp[5723]*kernel[0]+tmp[5724]*kernel[1]+tmp[5725]*kernel[2]+tmp[5823]*kernel[3]+tmp[5824]*kernel[4]+tmp[5825]*kernel[5]+tmp[5923]*kernel[6]+tmp[5924]*kernel[7]+tmp[5925]*kernel[8];
				ans[5825]<=tmp[5724]*kernel[0]+tmp[5725]*kernel[1]+tmp[5726]*kernel[2]+tmp[5824]*kernel[3]+tmp[5825]*kernel[4]+tmp[5826]*kernel[5]+tmp[5924]*kernel[6]+tmp[5925]*kernel[7]+tmp[5926]*kernel[8];
				ans[5826]<=tmp[5725]*kernel[0]+tmp[5726]*kernel[1]+tmp[5727]*kernel[2]+tmp[5825]*kernel[3]+tmp[5826]*kernel[4]+tmp[5827]*kernel[5]+tmp[5925]*kernel[6]+tmp[5926]*kernel[7]+tmp[5927]*kernel[8];
				ans[5827]<=tmp[5726]*kernel[0]+tmp[5727]*kernel[1]+tmp[5728]*kernel[2]+tmp[5826]*kernel[3]+tmp[5827]*kernel[4]+tmp[5828]*kernel[5]+tmp[5926]*kernel[6]+tmp[5927]*kernel[7]+tmp[5928]*kernel[8];
				ans[5828]<=tmp[5727]*kernel[0]+tmp[5728]*kernel[1]+tmp[5729]*kernel[2]+tmp[5827]*kernel[3]+tmp[5828]*kernel[4]+tmp[5829]*kernel[5]+tmp[5927]*kernel[6]+tmp[5928]*kernel[7]+tmp[5929]*kernel[8];
				ans[5829]<=tmp[5728]*kernel[0]+tmp[5729]*kernel[1]+tmp[5730]*kernel[2]+tmp[5828]*kernel[3]+tmp[5829]*kernel[4]+tmp[5830]*kernel[5]+tmp[5928]*kernel[6]+tmp[5929]*kernel[7]+tmp[5930]*kernel[8];
				ans[5830]<=tmp[5729]*kernel[0]+tmp[5730]*kernel[1]+tmp[5731]*kernel[2]+tmp[5829]*kernel[3]+tmp[5830]*kernel[4]+tmp[5831]*kernel[5]+tmp[5929]*kernel[6]+tmp[5930]*kernel[7]+tmp[5931]*kernel[8];
				ans[5831]<=tmp[5730]*kernel[0]+tmp[5731]*kernel[1]+tmp[5732]*kernel[2]+tmp[5830]*kernel[3]+tmp[5831]*kernel[4]+tmp[5832]*kernel[5]+tmp[5930]*kernel[6]+tmp[5931]*kernel[7]+tmp[5932]*kernel[8];
				ans[5832]<=tmp[5731]*kernel[0]+tmp[5732]*kernel[1]+tmp[5733]*kernel[2]+tmp[5831]*kernel[3]+tmp[5832]*kernel[4]+tmp[5833]*kernel[5]+tmp[5931]*kernel[6]+tmp[5932]*kernel[7]+tmp[5933]*kernel[8];
				ans[5833]<=tmp[5732]*kernel[0]+tmp[5733]*kernel[1]+tmp[5734]*kernel[2]+tmp[5832]*kernel[3]+tmp[5833]*kernel[4]+tmp[5834]*kernel[5]+tmp[5932]*kernel[6]+tmp[5933]*kernel[7]+tmp[5934]*kernel[8];
				ans[5834]<=tmp[5733]*kernel[0]+tmp[5734]*kernel[1]+tmp[5735]*kernel[2]+tmp[5833]*kernel[3]+tmp[5834]*kernel[4]+tmp[5835]*kernel[5]+tmp[5933]*kernel[6]+tmp[5934]*kernel[7]+tmp[5935]*kernel[8];
				ans[5835]<=tmp[5734]*kernel[0]+tmp[5735]*kernel[1]+tmp[5736]*kernel[2]+tmp[5834]*kernel[3]+tmp[5835]*kernel[4]+tmp[5836]*kernel[5]+tmp[5934]*kernel[6]+tmp[5935]*kernel[7]+tmp[5936]*kernel[8];
				ans[5836]<=tmp[5735]*kernel[0]+tmp[5736]*kernel[1]+tmp[5737]*kernel[2]+tmp[5835]*kernel[3]+tmp[5836]*kernel[4]+tmp[5837]*kernel[5]+tmp[5935]*kernel[6]+tmp[5936]*kernel[7]+tmp[5937]*kernel[8];
				ans[5837]<=tmp[5736]*kernel[0]+tmp[5737]*kernel[1]+tmp[5738]*kernel[2]+tmp[5836]*kernel[3]+tmp[5837]*kernel[4]+tmp[5838]*kernel[5]+tmp[5936]*kernel[6]+tmp[5937]*kernel[7]+tmp[5938]*kernel[8];
				ans[5838]<=tmp[5737]*kernel[0]+tmp[5738]*kernel[1]+tmp[5739]*kernel[2]+tmp[5837]*kernel[3]+tmp[5838]*kernel[4]+tmp[5839]*kernel[5]+tmp[5937]*kernel[6]+tmp[5938]*kernel[7]+tmp[5939]*kernel[8];
				ans[5839]<=tmp[5738]*kernel[0]+tmp[5739]*kernel[1]+tmp[5740]*kernel[2]+tmp[5838]*kernel[3]+tmp[5839]*kernel[4]+tmp[5840]*kernel[5]+tmp[5938]*kernel[6]+tmp[5939]*kernel[7]+tmp[5940]*kernel[8];
				ans[5840]<=tmp[5739]*kernel[0]+tmp[5740]*kernel[1]+tmp[5741]*kernel[2]+tmp[5839]*kernel[3]+tmp[5840]*kernel[4]+tmp[5841]*kernel[5]+tmp[5939]*kernel[6]+tmp[5940]*kernel[7]+tmp[5941]*kernel[8];
				ans[5841]<=tmp[5740]*kernel[0]+tmp[5741]*kernel[1]+tmp[5742]*kernel[2]+tmp[5840]*kernel[3]+tmp[5841]*kernel[4]+tmp[5842]*kernel[5]+tmp[5940]*kernel[6]+tmp[5941]*kernel[7]+tmp[5942]*kernel[8];
				ans[5842]<=tmp[5741]*kernel[0]+tmp[5742]*kernel[1]+tmp[5743]*kernel[2]+tmp[5841]*kernel[3]+tmp[5842]*kernel[4]+tmp[5843]*kernel[5]+tmp[5941]*kernel[6]+tmp[5942]*kernel[7]+tmp[5943]*kernel[8];
				ans[5843]<=tmp[5742]*kernel[0]+tmp[5743]*kernel[1]+tmp[5744]*kernel[2]+tmp[5842]*kernel[3]+tmp[5843]*kernel[4]+tmp[5844]*kernel[5]+tmp[5942]*kernel[6]+tmp[5943]*kernel[7]+tmp[5944]*kernel[8];
				ans[5844]<=tmp[5743]*kernel[0]+tmp[5744]*kernel[1]+tmp[5745]*kernel[2]+tmp[5843]*kernel[3]+tmp[5844]*kernel[4]+tmp[5845]*kernel[5]+tmp[5943]*kernel[6]+tmp[5944]*kernel[7]+tmp[5945]*kernel[8];
				ans[5845]<=tmp[5744]*kernel[0]+tmp[5745]*kernel[1]+tmp[5746]*kernel[2]+tmp[5844]*kernel[3]+tmp[5845]*kernel[4]+tmp[5846]*kernel[5]+tmp[5944]*kernel[6]+tmp[5945]*kernel[7]+tmp[5946]*kernel[8];
				ans[5846]<=tmp[5745]*kernel[0]+tmp[5746]*kernel[1]+tmp[5747]*kernel[2]+tmp[5845]*kernel[3]+tmp[5846]*kernel[4]+tmp[5847]*kernel[5]+tmp[5945]*kernel[6]+tmp[5946]*kernel[7]+tmp[5947]*kernel[8];
				ans[5847]<=tmp[5746]*kernel[0]+tmp[5747]*kernel[1]+tmp[5748]*kernel[2]+tmp[5846]*kernel[3]+tmp[5847]*kernel[4]+tmp[5848]*kernel[5]+tmp[5946]*kernel[6]+tmp[5947]*kernel[7]+tmp[5948]*kernel[8];
				ans[5848]<=tmp[5747]*kernel[0]+tmp[5748]*kernel[1]+tmp[5749]*kernel[2]+tmp[5847]*kernel[3]+tmp[5848]*kernel[4]+tmp[5849]*kernel[5]+tmp[5947]*kernel[6]+tmp[5948]*kernel[7]+tmp[5949]*kernel[8];
				ans[5849]<=tmp[5748]*kernel[0]+tmp[5749]*kernel[1]+tmp[5750]*kernel[2]+tmp[5848]*kernel[3]+tmp[5849]*kernel[4]+tmp[5850]*kernel[5]+tmp[5948]*kernel[6]+tmp[5949]*kernel[7]+tmp[5950]*kernel[8];
				ans[5850]<=tmp[5749]*kernel[0]+tmp[5750]*kernel[1]+tmp[5751]*kernel[2]+tmp[5849]*kernel[3]+tmp[5850]*kernel[4]+tmp[5851]*kernel[5]+tmp[5949]*kernel[6]+tmp[5950]*kernel[7]+tmp[5951]*kernel[8];
				ans[5851]<=tmp[5750]*kernel[0]+tmp[5751]*kernel[1]+tmp[5752]*kernel[2]+tmp[5850]*kernel[3]+tmp[5851]*kernel[4]+tmp[5852]*kernel[5]+tmp[5950]*kernel[6]+tmp[5951]*kernel[7]+tmp[5952]*kernel[8];
				ans[5852]<=tmp[5751]*kernel[0]+tmp[5752]*kernel[1]+tmp[5753]*kernel[2]+tmp[5851]*kernel[3]+tmp[5852]*kernel[4]+tmp[5853]*kernel[5]+tmp[5951]*kernel[6]+tmp[5952]*kernel[7]+tmp[5953]*kernel[8];
				ans[5853]<=tmp[5752]*kernel[0]+tmp[5753]*kernel[1]+tmp[5754]*kernel[2]+tmp[5852]*kernel[3]+tmp[5853]*kernel[4]+tmp[5854]*kernel[5]+tmp[5952]*kernel[6]+tmp[5953]*kernel[7]+tmp[5954]*kernel[8];
				ans[5854]<=tmp[5753]*kernel[0]+tmp[5754]*kernel[1]+tmp[5755]*kernel[2]+tmp[5853]*kernel[3]+tmp[5854]*kernel[4]+tmp[5855]*kernel[5]+tmp[5953]*kernel[6]+tmp[5954]*kernel[7]+tmp[5955]*kernel[8];
				ans[5855]<=tmp[5754]*kernel[0]+tmp[5755]*kernel[1]+tmp[5756]*kernel[2]+tmp[5854]*kernel[3]+tmp[5855]*kernel[4]+tmp[5856]*kernel[5]+tmp[5954]*kernel[6]+tmp[5955]*kernel[7]+tmp[5956]*kernel[8];
				ans[5856]<=tmp[5755]*kernel[0]+tmp[5756]*kernel[1]+tmp[5757]*kernel[2]+tmp[5855]*kernel[3]+tmp[5856]*kernel[4]+tmp[5857]*kernel[5]+tmp[5955]*kernel[6]+tmp[5956]*kernel[7]+tmp[5957]*kernel[8];
				ans[5857]<=tmp[5756]*kernel[0]+tmp[5757]*kernel[1]+tmp[5758]*kernel[2]+tmp[5856]*kernel[3]+tmp[5857]*kernel[4]+tmp[5858]*kernel[5]+tmp[5956]*kernel[6]+tmp[5957]*kernel[7]+tmp[5958]*kernel[8];
				ans[5858]<=tmp[5757]*kernel[0]+tmp[5758]*kernel[1]+tmp[5759]*kernel[2]+tmp[5857]*kernel[3]+tmp[5858]*kernel[4]+tmp[5859]*kernel[5]+tmp[5957]*kernel[6]+tmp[5958]*kernel[7]+tmp[5959]*kernel[8];
				ans[5859]<=tmp[5758]*kernel[0]+tmp[5759]*kernel[1]+tmp[5760]*kernel[2]+tmp[5858]*kernel[3]+tmp[5859]*kernel[4]+tmp[5860]*kernel[5]+tmp[5958]*kernel[6]+tmp[5959]*kernel[7]+tmp[5960]*kernel[8];
				ans[5860]<=tmp[5759]*kernel[0]+tmp[5760]*kernel[1]+tmp[5761]*kernel[2]+tmp[5859]*kernel[3]+tmp[5860]*kernel[4]+tmp[5861]*kernel[5]+tmp[5959]*kernel[6]+tmp[5960]*kernel[7]+tmp[5961]*kernel[8];
				ans[5861]<=tmp[5760]*kernel[0]+tmp[5761]*kernel[1]+tmp[5762]*kernel[2]+tmp[5860]*kernel[3]+tmp[5861]*kernel[4]+tmp[5862]*kernel[5]+tmp[5960]*kernel[6]+tmp[5961]*kernel[7]+tmp[5962]*kernel[8];
				ans[5862]<=tmp[5761]*kernel[0]+tmp[5762]*kernel[1]+tmp[5763]*kernel[2]+tmp[5861]*kernel[3]+tmp[5862]*kernel[4]+tmp[5863]*kernel[5]+tmp[5961]*kernel[6]+tmp[5962]*kernel[7]+tmp[5963]*kernel[8];
				ans[5863]<=tmp[5762]*kernel[0]+tmp[5763]*kernel[1]+tmp[5764]*kernel[2]+tmp[5862]*kernel[3]+tmp[5863]*kernel[4]+tmp[5864]*kernel[5]+tmp[5962]*kernel[6]+tmp[5963]*kernel[7]+tmp[5964]*kernel[8];
				ans[5864]<=tmp[5763]*kernel[0]+tmp[5764]*kernel[1]+tmp[5765]*kernel[2]+tmp[5863]*kernel[3]+tmp[5864]*kernel[4]+tmp[5865]*kernel[5]+tmp[5963]*kernel[6]+tmp[5964]*kernel[7]+tmp[5965]*kernel[8];
				ans[5865]<=tmp[5764]*kernel[0]+tmp[5765]*kernel[1]+tmp[5766]*kernel[2]+tmp[5864]*kernel[3]+tmp[5865]*kernel[4]+tmp[5866]*kernel[5]+tmp[5964]*kernel[6]+tmp[5965]*kernel[7]+tmp[5966]*kernel[8];
				ans[5866]<=tmp[5765]*kernel[0]+tmp[5766]*kernel[1]+tmp[5767]*kernel[2]+tmp[5865]*kernel[3]+tmp[5866]*kernel[4]+tmp[5867]*kernel[5]+tmp[5965]*kernel[6]+tmp[5966]*kernel[7]+tmp[5967]*kernel[8];
				ans[5867]<=tmp[5766]*kernel[0]+tmp[5767]*kernel[1]+tmp[5768]*kernel[2]+tmp[5866]*kernel[3]+tmp[5867]*kernel[4]+tmp[5868]*kernel[5]+tmp[5966]*kernel[6]+tmp[5967]*kernel[7]+tmp[5968]*kernel[8];
				ans[5868]<=tmp[5767]*kernel[0]+tmp[5768]*kernel[1]+tmp[5769]*kernel[2]+tmp[5867]*kernel[3]+tmp[5868]*kernel[4]+tmp[5869]*kernel[5]+tmp[5967]*kernel[6]+tmp[5968]*kernel[7]+tmp[5969]*kernel[8];
				ans[5869]<=tmp[5768]*kernel[0]+tmp[5769]*kernel[1]+tmp[5770]*kernel[2]+tmp[5868]*kernel[3]+tmp[5869]*kernel[4]+tmp[5870]*kernel[5]+tmp[5968]*kernel[6]+tmp[5969]*kernel[7]+tmp[5970]*kernel[8];
				ans[5870]<=tmp[5769]*kernel[0]+tmp[5770]*kernel[1]+tmp[5771]*kernel[2]+tmp[5869]*kernel[3]+tmp[5870]*kernel[4]+tmp[5871]*kernel[5]+tmp[5969]*kernel[6]+tmp[5970]*kernel[7]+tmp[5971]*kernel[8];
				ans[5871]<=tmp[5770]*kernel[0]+tmp[5771]*kernel[1]+tmp[5772]*kernel[2]+tmp[5870]*kernel[3]+tmp[5871]*kernel[4]+tmp[5872]*kernel[5]+tmp[5970]*kernel[6]+tmp[5971]*kernel[7]+tmp[5972]*kernel[8];
				ans[5872]<=tmp[5771]*kernel[0]+tmp[5772]*kernel[1]+tmp[5773]*kernel[2]+tmp[5871]*kernel[3]+tmp[5872]*kernel[4]+tmp[5873]*kernel[5]+tmp[5971]*kernel[6]+tmp[5972]*kernel[7]+tmp[5973]*kernel[8];
				ans[5873]<=tmp[5772]*kernel[0]+tmp[5773]*kernel[1]+tmp[5774]*kernel[2]+tmp[5872]*kernel[3]+tmp[5873]*kernel[4]+tmp[5874]*kernel[5]+tmp[5972]*kernel[6]+tmp[5973]*kernel[7]+tmp[5974]*kernel[8];
				ans[5874]<=tmp[5773]*kernel[0]+tmp[5774]*kernel[1]+tmp[5775]*kernel[2]+tmp[5873]*kernel[3]+tmp[5874]*kernel[4]+tmp[5875]*kernel[5]+tmp[5973]*kernel[6]+tmp[5974]*kernel[7]+tmp[5975]*kernel[8];
				ans[5875]<=tmp[5774]*kernel[0]+tmp[5775]*kernel[1]+tmp[5776]*kernel[2]+tmp[5874]*kernel[3]+tmp[5875]*kernel[4]+tmp[5876]*kernel[5]+tmp[5974]*kernel[6]+tmp[5975]*kernel[7]+tmp[5976]*kernel[8];
				ans[5876]<=tmp[5775]*kernel[0]+tmp[5776]*kernel[1]+tmp[5777]*kernel[2]+tmp[5875]*kernel[3]+tmp[5876]*kernel[4]+tmp[5877]*kernel[5]+tmp[5975]*kernel[6]+tmp[5976]*kernel[7]+tmp[5977]*kernel[8];
				ans[5877]<=tmp[5776]*kernel[0]+tmp[5777]*kernel[1]+tmp[5778]*kernel[2]+tmp[5876]*kernel[3]+tmp[5877]*kernel[4]+tmp[5878]*kernel[5]+tmp[5976]*kernel[6]+tmp[5977]*kernel[7]+tmp[5978]*kernel[8];
				ans[5878]<=tmp[5777]*kernel[0]+tmp[5778]*kernel[1]+tmp[5779]*kernel[2]+tmp[5877]*kernel[3]+tmp[5878]*kernel[4]+tmp[5879]*kernel[5]+tmp[5977]*kernel[6]+tmp[5978]*kernel[7]+tmp[5979]*kernel[8];
				ans[5879]<=tmp[5778]*kernel[0]+tmp[5779]*kernel[1]+tmp[5780]*kernel[2]+tmp[5878]*kernel[3]+tmp[5879]*kernel[4]+tmp[5880]*kernel[5]+tmp[5978]*kernel[6]+tmp[5979]*kernel[7]+tmp[5980]*kernel[8];
				ans[5880]<=tmp[5779]*kernel[0]+tmp[5780]*kernel[1]+tmp[5781]*kernel[2]+tmp[5879]*kernel[3]+tmp[5880]*kernel[4]+tmp[5881]*kernel[5]+tmp[5979]*kernel[6]+tmp[5980]*kernel[7]+tmp[5981]*kernel[8];
				ans[5881]<=tmp[5780]*kernel[0]+tmp[5781]*kernel[1]+tmp[5782]*kernel[2]+tmp[5880]*kernel[3]+tmp[5881]*kernel[4]+tmp[5882]*kernel[5]+tmp[5980]*kernel[6]+tmp[5981]*kernel[7]+tmp[5982]*kernel[8];
				ans[5882]<=tmp[5781]*kernel[0]+tmp[5782]*kernel[1]+tmp[5783]*kernel[2]+tmp[5881]*kernel[3]+tmp[5882]*kernel[4]+tmp[5883]*kernel[5]+tmp[5981]*kernel[6]+tmp[5982]*kernel[7]+tmp[5983]*kernel[8];
				ans[5883]<=tmp[5782]*kernel[0]+tmp[5783]*kernel[1]+tmp[5784]*kernel[2]+tmp[5882]*kernel[3]+tmp[5883]*kernel[4]+tmp[5884]*kernel[5]+tmp[5982]*kernel[6]+tmp[5983]*kernel[7]+tmp[5984]*kernel[8];
				ans[5884]<=tmp[5783]*kernel[0]+tmp[5784]*kernel[1]+tmp[5785]*kernel[2]+tmp[5883]*kernel[3]+tmp[5884]*kernel[4]+tmp[5885]*kernel[5]+tmp[5983]*kernel[6]+tmp[5984]*kernel[7]+tmp[5985]*kernel[8];
				ans[5885]<=tmp[5784]*kernel[0]+tmp[5785]*kernel[1]+tmp[5786]*kernel[2]+tmp[5884]*kernel[3]+tmp[5885]*kernel[4]+tmp[5886]*kernel[5]+tmp[5984]*kernel[6]+tmp[5985]*kernel[7]+tmp[5986]*kernel[8];
				ans[5886]<=tmp[5785]*kernel[0]+tmp[5786]*kernel[1]+tmp[5787]*kernel[2]+tmp[5885]*kernel[3]+tmp[5886]*kernel[4]+tmp[5887]*kernel[5]+tmp[5985]*kernel[6]+tmp[5986]*kernel[7]+tmp[5987]*kernel[8];
				ans[5887]<=tmp[5786]*kernel[0]+tmp[5787]*kernel[1]+tmp[5788]*kernel[2]+tmp[5886]*kernel[3]+tmp[5887]*kernel[4]+tmp[5888]*kernel[5]+tmp[5986]*kernel[6]+tmp[5987]*kernel[7]+tmp[5988]*kernel[8];
				ans[5888]<=tmp[5787]*kernel[0]+tmp[5788]*kernel[1]+tmp[5789]*kernel[2]+tmp[5887]*kernel[3]+tmp[5888]*kernel[4]+tmp[5889]*kernel[5]+tmp[5987]*kernel[6]+tmp[5988]*kernel[7]+tmp[5989]*kernel[8];
				ans[5889]<=tmp[5788]*kernel[0]+tmp[5789]*kernel[1]+tmp[5790]*kernel[2]+tmp[5888]*kernel[3]+tmp[5889]*kernel[4]+tmp[5890]*kernel[5]+tmp[5988]*kernel[6]+tmp[5989]*kernel[7]+tmp[5990]*kernel[8];
				ans[5890]<=tmp[5789]*kernel[0]+tmp[5790]*kernel[1]+tmp[5791]*kernel[2]+tmp[5889]*kernel[3]+tmp[5890]*kernel[4]+tmp[5891]*kernel[5]+tmp[5989]*kernel[6]+tmp[5990]*kernel[7]+tmp[5991]*kernel[8];
				ans[5891]<=tmp[5790]*kernel[0]+tmp[5791]*kernel[1]+tmp[5792]*kernel[2]+tmp[5890]*kernel[3]+tmp[5891]*kernel[4]+tmp[5892]*kernel[5]+tmp[5990]*kernel[6]+tmp[5991]*kernel[7]+tmp[5992]*kernel[8];
				ans[5892]<=tmp[5791]*kernel[0]+tmp[5792]*kernel[1]+tmp[5793]*kernel[2]+tmp[5891]*kernel[3]+tmp[5892]*kernel[4]+tmp[5893]*kernel[5]+tmp[5991]*kernel[6]+tmp[5992]*kernel[7]+tmp[5993]*kernel[8];
				ans[5893]<=tmp[5792]*kernel[0]+tmp[5793]*kernel[1]+tmp[5794]*kernel[2]+tmp[5892]*kernel[3]+tmp[5893]*kernel[4]+tmp[5894]*kernel[5]+tmp[5992]*kernel[6]+tmp[5993]*kernel[7]+tmp[5994]*kernel[8];
				ans[5894]<=tmp[5793]*kernel[0]+tmp[5794]*kernel[1]+tmp[5795]*kernel[2]+tmp[5893]*kernel[3]+tmp[5894]*kernel[4]+tmp[5895]*kernel[5]+tmp[5993]*kernel[6]+tmp[5994]*kernel[7]+tmp[5995]*kernel[8];
				ans[5895]<=tmp[5794]*kernel[0]+tmp[5795]*kernel[1]+tmp[5796]*kernel[2]+tmp[5894]*kernel[3]+tmp[5895]*kernel[4]+tmp[5896]*kernel[5]+tmp[5994]*kernel[6]+tmp[5995]*kernel[7]+tmp[5996]*kernel[8];
				ans[5896]<=tmp[5795]*kernel[0]+tmp[5796]*kernel[1]+tmp[5797]*kernel[2]+tmp[5895]*kernel[3]+tmp[5896]*kernel[4]+tmp[5897]*kernel[5]+tmp[5995]*kernel[6]+tmp[5996]*kernel[7]+tmp[5997]*kernel[8];
				ans[5897]<=tmp[5796]*kernel[0]+tmp[5797]*kernel[1]+tmp[5798]*kernel[2]+tmp[5896]*kernel[3]+tmp[5897]*kernel[4]+tmp[5898]*kernel[5]+tmp[5996]*kernel[6]+tmp[5997]*kernel[7]+tmp[5998]*kernel[8];
				ans[5898]<=tmp[5797]*kernel[0]+tmp[5798]*kernel[1]+tmp[5799]*kernel[2]+tmp[5897]*kernel[3]+tmp[5898]*kernel[4]+tmp[5899]*kernel[5]+tmp[5997]*kernel[6]+tmp[5998]*kernel[7]+tmp[5999]*kernel[8];
				ans[5899]<=tmp[5798]*kernel[0]+tmp[5799]*kernel[1]+tmp[5898]*kernel[3]+tmp[5899]*kernel[4]+tmp[5998]*kernel[6]+tmp[5999]*kernel[7];
				ans[5900]<=tmp[5800]*kernel[1]+tmp[5801]*kernel[2]+tmp[5900]*kernel[4]+tmp[5901]*kernel[5]+tmp[6000]*kernel[7]+tmp[6001]*kernel[8];
				ans[5901]<=tmp[5800]*kernel[0]+tmp[5801]*kernel[1]+tmp[5802]*kernel[2]+tmp[5900]*kernel[3]+tmp[5901]*kernel[4]+tmp[5902]*kernel[5]+tmp[6000]*kernel[6]+tmp[6001]*kernel[7]+tmp[6002]*kernel[8];
				ans[5902]<=tmp[5801]*kernel[0]+tmp[5802]*kernel[1]+tmp[5803]*kernel[2]+tmp[5901]*kernel[3]+tmp[5902]*kernel[4]+tmp[5903]*kernel[5]+tmp[6001]*kernel[6]+tmp[6002]*kernel[7]+tmp[6003]*kernel[8];
				ans[5903]<=tmp[5802]*kernel[0]+tmp[5803]*kernel[1]+tmp[5804]*kernel[2]+tmp[5902]*kernel[3]+tmp[5903]*kernel[4]+tmp[5904]*kernel[5]+tmp[6002]*kernel[6]+tmp[6003]*kernel[7]+tmp[6004]*kernel[8];
				ans[5904]<=tmp[5803]*kernel[0]+tmp[5804]*kernel[1]+tmp[5805]*kernel[2]+tmp[5903]*kernel[3]+tmp[5904]*kernel[4]+tmp[5905]*kernel[5]+tmp[6003]*kernel[6]+tmp[6004]*kernel[7]+tmp[6005]*kernel[8];
				ans[5905]<=tmp[5804]*kernel[0]+tmp[5805]*kernel[1]+tmp[5806]*kernel[2]+tmp[5904]*kernel[3]+tmp[5905]*kernel[4]+tmp[5906]*kernel[5]+tmp[6004]*kernel[6]+tmp[6005]*kernel[7]+tmp[6006]*kernel[8];
				ans[5906]<=tmp[5805]*kernel[0]+tmp[5806]*kernel[1]+tmp[5807]*kernel[2]+tmp[5905]*kernel[3]+tmp[5906]*kernel[4]+tmp[5907]*kernel[5]+tmp[6005]*kernel[6]+tmp[6006]*kernel[7]+tmp[6007]*kernel[8];
				ans[5907]<=tmp[5806]*kernel[0]+tmp[5807]*kernel[1]+tmp[5808]*kernel[2]+tmp[5906]*kernel[3]+tmp[5907]*kernel[4]+tmp[5908]*kernel[5]+tmp[6006]*kernel[6]+tmp[6007]*kernel[7]+tmp[6008]*kernel[8];
				ans[5908]<=tmp[5807]*kernel[0]+tmp[5808]*kernel[1]+tmp[5809]*kernel[2]+tmp[5907]*kernel[3]+tmp[5908]*kernel[4]+tmp[5909]*kernel[5]+tmp[6007]*kernel[6]+tmp[6008]*kernel[7]+tmp[6009]*kernel[8];
				ans[5909]<=tmp[5808]*kernel[0]+tmp[5809]*kernel[1]+tmp[5810]*kernel[2]+tmp[5908]*kernel[3]+tmp[5909]*kernel[4]+tmp[5910]*kernel[5]+tmp[6008]*kernel[6]+tmp[6009]*kernel[7]+tmp[6010]*kernel[8];
				ans[5910]<=tmp[5809]*kernel[0]+tmp[5810]*kernel[1]+tmp[5811]*kernel[2]+tmp[5909]*kernel[3]+tmp[5910]*kernel[4]+tmp[5911]*kernel[5]+tmp[6009]*kernel[6]+tmp[6010]*kernel[7]+tmp[6011]*kernel[8];
				ans[5911]<=tmp[5810]*kernel[0]+tmp[5811]*kernel[1]+tmp[5812]*kernel[2]+tmp[5910]*kernel[3]+tmp[5911]*kernel[4]+tmp[5912]*kernel[5]+tmp[6010]*kernel[6]+tmp[6011]*kernel[7]+tmp[6012]*kernel[8];
				ans[5912]<=tmp[5811]*kernel[0]+tmp[5812]*kernel[1]+tmp[5813]*kernel[2]+tmp[5911]*kernel[3]+tmp[5912]*kernel[4]+tmp[5913]*kernel[5]+tmp[6011]*kernel[6]+tmp[6012]*kernel[7]+tmp[6013]*kernel[8];
				ans[5913]<=tmp[5812]*kernel[0]+tmp[5813]*kernel[1]+tmp[5814]*kernel[2]+tmp[5912]*kernel[3]+tmp[5913]*kernel[4]+tmp[5914]*kernel[5]+tmp[6012]*kernel[6]+tmp[6013]*kernel[7]+tmp[6014]*kernel[8];
				ans[5914]<=tmp[5813]*kernel[0]+tmp[5814]*kernel[1]+tmp[5815]*kernel[2]+tmp[5913]*kernel[3]+tmp[5914]*kernel[4]+tmp[5915]*kernel[5]+tmp[6013]*kernel[6]+tmp[6014]*kernel[7]+tmp[6015]*kernel[8];
				ans[5915]<=tmp[5814]*kernel[0]+tmp[5815]*kernel[1]+tmp[5816]*kernel[2]+tmp[5914]*kernel[3]+tmp[5915]*kernel[4]+tmp[5916]*kernel[5]+tmp[6014]*kernel[6]+tmp[6015]*kernel[7]+tmp[6016]*kernel[8];
				ans[5916]<=tmp[5815]*kernel[0]+tmp[5816]*kernel[1]+tmp[5817]*kernel[2]+tmp[5915]*kernel[3]+tmp[5916]*kernel[4]+tmp[5917]*kernel[5]+tmp[6015]*kernel[6]+tmp[6016]*kernel[7]+tmp[6017]*kernel[8];
				ans[5917]<=tmp[5816]*kernel[0]+tmp[5817]*kernel[1]+tmp[5818]*kernel[2]+tmp[5916]*kernel[3]+tmp[5917]*kernel[4]+tmp[5918]*kernel[5]+tmp[6016]*kernel[6]+tmp[6017]*kernel[7]+tmp[6018]*kernel[8];
				ans[5918]<=tmp[5817]*kernel[0]+tmp[5818]*kernel[1]+tmp[5819]*kernel[2]+tmp[5917]*kernel[3]+tmp[5918]*kernel[4]+tmp[5919]*kernel[5]+tmp[6017]*kernel[6]+tmp[6018]*kernel[7]+tmp[6019]*kernel[8];
				ans[5919]<=tmp[5818]*kernel[0]+tmp[5819]*kernel[1]+tmp[5820]*kernel[2]+tmp[5918]*kernel[3]+tmp[5919]*kernel[4]+tmp[5920]*kernel[5]+tmp[6018]*kernel[6]+tmp[6019]*kernel[7]+tmp[6020]*kernel[8];
				ans[5920]<=tmp[5819]*kernel[0]+tmp[5820]*kernel[1]+tmp[5821]*kernel[2]+tmp[5919]*kernel[3]+tmp[5920]*kernel[4]+tmp[5921]*kernel[5]+tmp[6019]*kernel[6]+tmp[6020]*kernel[7]+tmp[6021]*kernel[8];
				ans[5921]<=tmp[5820]*kernel[0]+tmp[5821]*kernel[1]+tmp[5822]*kernel[2]+tmp[5920]*kernel[3]+tmp[5921]*kernel[4]+tmp[5922]*kernel[5]+tmp[6020]*kernel[6]+tmp[6021]*kernel[7]+tmp[6022]*kernel[8];
				ans[5922]<=tmp[5821]*kernel[0]+tmp[5822]*kernel[1]+tmp[5823]*kernel[2]+tmp[5921]*kernel[3]+tmp[5922]*kernel[4]+tmp[5923]*kernel[5]+tmp[6021]*kernel[6]+tmp[6022]*kernel[7]+tmp[6023]*kernel[8];
				ans[5923]<=tmp[5822]*kernel[0]+tmp[5823]*kernel[1]+tmp[5824]*kernel[2]+tmp[5922]*kernel[3]+tmp[5923]*kernel[4]+tmp[5924]*kernel[5]+tmp[6022]*kernel[6]+tmp[6023]*kernel[7]+tmp[6024]*kernel[8];
				ans[5924]<=tmp[5823]*kernel[0]+tmp[5824]*kernel[1]+tmp[5825]*kernel[2]+tmp[5923]*kernel[3]+tmp[5924]*kernel[4]+tmp[5925]*kernel[5]+tmp[6023]*kernel[6]+tmp[6024]*kernel[7]+tmp[6025]*kernel[8];
				ans[5925]<=tmp[5824]*kernel[0]+tmp[5825]*kernel[1]+tmp[5826]*kernel[2]+tmp[5924]*kernel[3]+tmp[5925]*kernel[4]+tmp[5926]*kernel[5]+tmp[6024]*kernel[6]+tmp[6025]*kernel[7]+tmp[6026]*kernel[8];
				ans[5926]<=tmp[5825]*kernel[0]+tmp[5826]*kernel[1]+tmp[5827]*kernel[2]+tmp[5925]*kernel[3]+tmp[5926]*kernel[4]+tmp[5927]*kernel[5]+tmp[6025]*kernel[6]+tmp[6026]*kernel[7]+tmp[6027]*kernel[8];
				ans[5927]<=tmp[5826]*kernel[0]+tmp[5827]*kernel[1]+tmp[5828]*kernel[2]+tmp[5926]*kernel[3]+tmp[5927]*kernel[4]+tmp[5928]*kernel[5]+tmp[6026]*kernel[6]+tmp[6027]*kernel[7]+tmp[6028]*kernel[8];
				ans[5928]<=tmp[5827]*kernel[0]+tmp[5828]*kernel[1]+tmp[5829]*kernel[2]+tmp[5927]*kernel[3]+tmp[5928]*kernel[4]+tmp[5929]*kernel[5]+tmp[6027]*kernel[6]+tmp[6028]*kernel[7]+tmp[6029]*kernel[8];
				ans[5929]<=tmp[5828]*kernel[0]+tmp[5829]*kernel[1]+tmp[5830]*kernel[2]+tmp[5928]*kernel[3]+tmp[5929]*kernel[4]+tmp[5930]*kernel[5]+tmp[6028]*kernel[6]+tmp[6029]*kernel[7]+tmp[6030]*kernel[8];
				ans[5930]<=tmp[5829]*kernel[0]+tmp[5830]*kernel[1]+tmp[5831]*kernel[2]+tmp[5929]*kernel[3]+tmp[5930]*kernel[4]+tmp[5931]*kernel[5]+tmp[6029]*kernel[6]+tmp[6030]*kernel[7]+tmp[6031]*kernel[8];
				ans[5931]<=tmp[5830]*kernel[0]+tmp[5831]*kernel[1]+tmp[5832]*kernel[2]+tmp[5930]*kernel[3]+tmp[5931]*kernel[4]+tmp[5932]*kernel[5]+tmp[6030]*kernel[6]+tmp[6031]*kernel[7]+tmp[6032]*kernel[8];
				ans[5932]<=tmp[5831]*kernel[0]+tmp[5832]*kernel[1]+tmp[5833]*kernel[2]+tmp[5931]*kernel[3]+tmp[5932]*kernel[4]+tmp[5933]*kernel[5]+tmp[6031]*kernel[6]+tmp[6032]*kernel[7]+tmp[6033]*kernel[8];
				ans[5933]<=tmp[5832]*kernel[0]+tmp[5833]*kernel[1]+tmp[5834]*kernel[2]+tmp[5932]*kernel[3]+tmp[5933]*kernel[4]+tmp[5934]*kernel[5]+tmp[6032]*kernel[6]+tmp[6033]*kernel[7]+tmp[6034]*kernel[8];
				ans[5934]<=tmp[5833]*kernel[0]+tmp[5834]*kernel[1]+tmp[5835]*kernel[2]+tmp[5933]*kernel[3]+tmp[5934]*kernel[4]+tmp[5935]*kernel[5]+tmp[6033]*kernel[6]+tmp[6034]*kernel[7]+tmp[6035]*kernel[8];
				ans[5935]<=tmp[5834]*kernel[0]+tmp[5835]*kernel[1]+tmp[5836]*kernel[2]+tmp[5934]*kernel[3]+tmp[5935]*kernel[4]+tmp[5936]*kernel[5]+tmp[6034]*kernel[6]+tmp[6035]*kernel[7]+tmp[6036]*kernel[8];
				ans[5936]<=tmp[5835]*kernel[0]+tmp[5836]*kernel[1]+tmp[5837]*kernel[2]+tmp[5935]*kernel[3]+tmp[5936]*kernel[4]+tmp[5937]*kernel[5]+tmp[6035]*kernel[6]+tmp[6036]*kernel[7]+tmp[6037]*kernel[8];
				ans[5937]<=tmp[5836]*kernel[0]+tmp[5837]*kernel[1]+tmp[5838]*kernel[2]+tmp[5936]*kernel[3]+tmp[5937]*kernel[4]+tmp[5938]*kernel[5]+tmp[6036]*kernel[6]+tmp[6037]*kernel[7]+tmp[6038]*kernel[8];
				ans[5938]<=tmp[5837]*kernel[0]+tmp[5838]*kernel[1]+tmp[5839]*kernel[2]+tmp[5937]*kernel[3]+tmp[5938]*kernel[4]+tmp[5939]*kernel[5]+tmp[6037]*kernel[6]+tmp[6038]*kernel[7]+tmp[6039]*kernel[8];
				ans[5939]<=tmp[5838]*kernel[0]+tmp[5839]*kernel[1]+tmp[5840]*kernel[2]+tmp[5938]*kernel[3]+tmp[5939]*kernel[4]+tmp[5940]*kernel[5]+tmp[6038]*kernel[6]+tmp[6039]*kernel[7]+tmp[6040]*kernel[8];
				ans[5940]<=tmp[5839]*kernel[0]+tmp[5840]*kernel[1]+tmp[5841]*kernel[2]+tmp[5939]*kernel[3]+tmp[5940]*kernel[4]+tmp[5941]*kernel[5]+tmp[6039]*kernel[6]+tmp[6040]*kernel[7]+tmp[6041]*kernel[8];
				ans[5941]<=tmp[5840]*kernel[0]+tmp[5841]*kernel[1]+tmp[5842]*kernel[2]+tmp[5940]*kernel[3]+tmp[5941]*kernel[4]+tmp[5942]*kernel[5]+tmp[6040]*kernel[6]+tmp[6041]*kernel[7]+tmp[6042]*kernel[8];
				ans[5942]<=tmp[5841]*kernel[0]+tmp[5842]*kernel[1]+tmp[5843]*kernel[2]+tmp[5941]*kernel[3]+tmp[5942]*kernel[4]+tmp[5943]*kernel[5]+tmp[6041]*kernel[6]+tmp[6042]*kernel[7]+tmp[6043]*kernel[8];
				ans[5943]<=tmp[5842]*kernel[0]+tmp[5843]*kernel[1]+tmp[5844]*kernel[2]+tmp[5942]*kernel[3]+tmp[5943]*kernel[4]+tmp[5944]*kernel[5]+tmp[6042]*kernel[6]+tmp[6043]*kernel[7]+tmp[6044]*kernel[8];
				ans[5944]<=tmp[5843]*kernel[0]+tmp[5844]*kernel[1]+tmp[5845]*kernel[2]+tmp[5943]*kernel[3]+tmp[5944]*kernel[4]+tmp[5945]*kernel[5]+tmp[6043]*kernel[6]+tmp[6044]*kernel[7]+tmp[6045]*kernel[8];
				ans[5945]<=tmp[5844]*kernel[0]+tmp[5845]*kernel[1]+tmp[5846]*kernel[2]+tmp[5944]*kernel[3]+tmp[5945]*kernel[4]+tmp[5946]*kernel[5]+tmp[6044]*kernel[6]+tmp[6045]*kernel[7]+tmp[6046]*kernel[8];
				ans[5946]<=tmp[5845]*kernel[0]+tmp[5846]*kernel[1]+tmp[5847]*kernel[2]+tmp[5945]*kernel[3]+tmp[5946]*kernel[4]+tmp[5947]*kernel[5]+tmp[6045]*kernel[6]+tmp[6046]*kernel[7]+tmp[6047]*kernel[8];
				ans[5947]<=tmp[5846]*kernel[0]+tmp[5847]*kernel[1]+tmp[5848]*kernel[2]+tmp[5946]*kernel[3]+tmp[5947]*kernel[4]+tmp[5948]*kernel[5]+tmp[6046]*kernel[6]+tmp[6047]*kernel[7]+tmp[6048]*kernel[8];
				ans[5948]<=tmp[5847]*kernel[0]+tmp[5848]*kernel[1]+tmp[5849]*kernel[2]+tmp[5947]*kernel[3]+tmp[5948]*kernel[4]+tmp[5949]*kernel[5]+tmp[6047]*kernel[6]+tmp[6048]*kernel[7]+tmp[6049]*kernel[8];
				ans[5949]<=tmp[5848]*kernel[0]+tmp[5849]*kernel[1]+tmp[5850]*kernel[2]+tmp[5948]*kernel[3]+tmp[5949]*kernel[4]+tmp[5950]*kernel[5]+tmp[6048]*kernel[6]+tmp[6049]*kernel[7]+tmp[6050]*kernel[8];
				ans[5950]<=tmp[5849]*kernel[0]+tmp[5850]*kernel[1]+tmp[5851]*kernel[2]+tmp[5949]*kernel[3]+tmp[5950]*kernel[4]+tmp[5951]*kernel[5]+tmp[6049]*kernel[6]+tmp[6050]*kernel[7]+tmp[6051]*kernel[8];
				ans[5951]<=tmp[5850]*kernel[0]+tmp[5851]*kernel[1]+tmp[5852]*kernel[2]+tmp[5950]*kernel[3]+tmp[5951]*kernel[4]+tmp[5952]*kernel[5]+tmp[6050]*kernel[6]+tmp[6051]*kernel[7]+tmp[6052]*kernel[8];
				ans[5952]<=tmp[5851]*kernel[0]+tmp[5852]*kernel[1]+tmp[5853]*kernel[2]+tmp[5951]*kernel[3]+tmp[5952]*kernel[4]+tmp[5953]*kernel[5]+tmp[6051]*kernel[6]+tmp[6052]*kernel[7]+tmp[6053]*kernel[8];
				ans[5953]<=tmp[5852]*kernel[0]+tmp[5853]*kernel[1]+tmp[5854]*kernel[2]+tmp[5952]*kernel[3]+tmp[5953]*kernel[4]+tmp[5954]*kernel[5]+tmp[6052]*kernel[6]+tmp[6053]*kernel[7]+tmp[6054]*kernel[8];
				ans[5954]<=tmp[5853]*kernel[0]+tmp[5854]*kernel[1]+tmp[5855]*kernel[2]+tmp[5953]*kernel[3]+tmp[5954]*kernel[4]+tmp[5955]*kernel[5]+tmp[6053]*kernel[6]+tmp[6054]*kernel[7]+tmp[6055]*kernel[8];
				ans[5955]<=tmp[5854]*kernel[0]+tmp[5855]*kernel[1]+tmp[5856]*kernel[2]+tmp[5954]*kernel[3]+tmp[5955]*kernel[4]+tmp[5956]*kernel[5]+tmp[6054]*kernel[6]+tmp[6055]*kernel[7]+tmp[6056]*kernel[8];
				ans[5956]<=tmp[5855]*kernel[0]+tmp[5856]*kernel[1]+tmp[5857]*kernel[2]+tmp[5955]*kernel[3]+tmp[5956]*kernel[4]+tmp[5957]*kernel[5]+tmp[6055]*kernel[6]+tmp[6056]*kernel[7]+tmp[6057]*kernel[8];
				ans[5957]<=tmp[5856]*kernel[0]+tmp[5857]*kernel[1]+tmp[5858]*kernel[2]+tmp[5956]*kernel[3]+tmp[5957]*kernel[4]+tmp[5958]*kernel[5]+tmp[6056]*kernel[6]+tmp[6057]*kernel[7]+tmp[6058]*kernel[8];
				ans[5958]<=tmp[5857]*kernel[0]+tmp[5858]*kernel[1]+tmp[5859]*kernel[2]+tmp[5957]*kernel[3]+tmp[5958]*kernel[4]+tmp[5959]*kernel[5]+tmp[6057]*kernel[6]+tmp[6058]*kernel[7]+tmp[6059]*kernel[8];
				ans[5959]<=tmp[5858]*kernel[0]+tmp[5859]*kernel[1]+tmp[5860]*kernel[2]+tmp[5958]*kernel[3]+tmp[5959]*kernel[4]+tmp[5960]*kernel[5]+tmp[6058]*kernel[6]+tmp[6059]*kernel[7]+tmp[6060]*kernel[8];
				ans[5960]<=tmp[5859]*kernel[0]+tmp[5860]*kernel[1]+tmp[5861]*kernel[2]+tmp[5959]*kernel[3]+tmp[5960]*kernel[4]+tmp[5961]*kernel[5]+tmp[6059]*kernel[6]+tmp[6060]*kernel[7]+tmp[6061]*kernel[8];
				ans[5961]<=tmp[5860]*kernel[0]+tmp[5861]*kernel[1]+tmp[5862]*kernel[2]+tmp[5960]*kernel[3]+tmp[5961]*kernel[4]+tmp[5962]*kernel[5]+tmp[6060]*kernel[6]+tmp[6061]*kernel[7]+tmp[6062]*kernel[8];
				ans[5962]<=tmp[5861]*kernel[0]+tmp[5862]*kernel[1]+tmp[5863]*kernel[2]+tmp[5961]*kernel[3]+tmp[5962]*kernel[4]+tmp[5963]*kernel[5]+tmp[6061]*kernel[6]+tmp[6062]*kernel[7]+tmp[6063]*kernel[8];
				ans[5963]<=tmp[5862]*kernel[0]+tmp[5863]*kernel[1]+tmp[5864]*kernel[2]+tmp[5962]*kernel[3]+tmp[5963]*kernel[4]+tmp[5964]*kernel[5]+tmp[6062]*kernel[6]+tmp[6063]*kernel[7]+tmp[6064]*kernel[8];
				ans[5964]<=tmp[5863]*kernel[0]+tmp[5864]*kernel[1]+tmp[5865]*kernel[2]+tmp[5963]*kernel[3]+tmp[5964]*kernel[4]+tmp[5965]*kernel[5]+tmp[6063]*kernel[6]+tmp[6064]*kernel[7]+tmp[6065]*kernel[8];
				ans[5965]<=tmp[5864]*kernel[0]+tmp[5865]*kernel[1]+tmp[5866]*kernel[2]+tmp[5964]*kernel[3]+tmp[5965]*kernel[4]+tmp[5966]*kernel[5]+tmp[6064]*kernel[6]+tmp[6065]*kernel[7]+tmp[6066]*kernel[8];
				ans[5966]<=tmp[5865]*kernel[0]+tmp[5866]*kernel[1]+tmp[5867]*kernel[2]+tmp[5965]*kernel[3]+tmp[5966]*kernel[4]+tmp[5967]*kernel[5]+tmp[6065]*kernel[6]+tmp[6066]*kernel[7]+tmp[6067]*kernel[8];
				ans[5967]<=tmp[5866]*kernel[0]+tmp[5867]*kernel[1]+tmp[5868]*kernel[2]+tmp[5966]*kernel[3]+tmp[5967]*kernel[4]+tmp[5968]*kernel[5]+tmp[6066]*kernel[6]+tmp[6067]*kernel[7]+tmp[6068]*kernel[8];
				ans[5968]<=tmp[5867]*kernel[0]+tmp[5868]*kernel[1]+tmp[5869]*kernel[2]+tmp[5967]*kernel[3]+tmp[5968]*kernel[4]+tmp[5969]*kernel[5]+tmp[6067]*kernel[6]+tmp[6068]*kernel[7]+tmp[6069]*kernel[8];
				ans[5969]<=tmp[5868]*kernel[0]+tmp[5869]*kernel[1]+tmp[5870]*kernel[2]+tmp[5968]*kernel[3]+tmp[5969]*kernel[4]+tmp[5970]*kernel[5]+tmp[6068]*kernel[6]+tmp[6069]*kernel[7]+tmp[6070]*kernel[8];
				ans[5970]<=tmp[5869]*kernel[0]+tmp[5870]*kernel[1]+tmp[5871]*kernel[2]+tmp[5969]*kernel[3]+tmp[5970]*kernel[4]+tmp[5971]*kernel[5]+tmp[6069]*kernel[6]+tmp[6070]*kernel[7]+tmp[6071]*kernel[8];
				ans[5971]<=tmp[5870]*kernel[0]+tmp[5871]*kernel[1]+tmp[5872]*kernel[2]+tmp[5970]*kernel[3]+tmp[5971]*kernel[4]+tmp[5972]*kernel[5]+tmp[6070]*kernel[6]+tmp[6071]*kernel[7]+tmp[6072]*kernel[8];
				ans[5972]<=tmp[5871]*kernel[0]+tmp[5872]*kernel[1]+tmp[5873]*kernel[2]+tmp[5971]*kernel[3]+tmp[5972]*kernel[4]+tmp[5973]*kernel[5]+tmp[6071]*kernel[6]+tmp[6072]*kernel[7]+tmp[6073]*kernel[8];
				ans[5973]<=tmp[5872]*kernel[0]+tmp[5873]*kernel[1]+tmp[5874]*kernel[2]+tmp[5972]*kernel[3]+tmp[5973]*kernel[4]+tmp[5974]*kernel[5]+tmp[6072]*kernel[6]+tmp[6073]*kernel[7]+tmp[6074]*kernel[8];
				ans[5974]<=tmp[5873]*kernel[0]+tmp[5874]*kernel[1]+tmp[5875]*kernel[2]+tmp[5973]*kernel[3]+tmp[5974]*kernel[4]+tmp[5975]*kernel[5]+tmp[6073]*kernel[6]+tmp[6074]*kernel[7]+tmp[6075]*kernel[8];
				ans[5975]<=tmp[5874]*kernel[0]+tmp[5875]*kernel[1]+tmp[5876]*kernel[2]+tmp[5974]*kernel[3]+tmp[5975]*kernel[4]+tmp[5976]*kernel[5]+tmp[6074]*kernel[6]+tmp[6075]*kernel[7]+tmp[6076]*kernel[8];
				ans[5976]<=tmp[5875]*kernel[0]+tmp[5876]*kernel[1]+tmp[5877]*kernel[2]+tmp[5975]*kernel[3]+tmp[5976]*kernel[4]+tmp[5977]*kernel[5]+tmp[6075]*kernel[6]+tmp[6076]*kernel[7]+tmp[6077]*kernel[8];
				ans[5977]<=tmp[5876]*kernel[0]+tmp[5877]*kernel[1]+tmp[5878]*kernel[2]+tmp[5976]*kernel[3]+tmp[5977]*kernel[4]+tmp[5978]*kernel[5]+tmp[6076]*kernel[6]+tmp[6077]*kernel[7]+tmp[6078]*kernel[8];
				ans[5978]<=tmp[5877]*kernel[0]+tmp[5878]*kernel[1]+tmp[5879]*kernel[2]+tmp[5977]*kernel[3]+tmp[5978]*kernel[4]+tmp[5979]*kernel[5]+tmp[6077]*kernel[6]+tmp[6078]*kernel[7]+tmp[6079]*kernel[8];
				ans[5979]<=tmp[5878]*kernel[0]+tmp[5879]*kernel[1]+tmp[5880]*kernel[2]+tmp[5978]*kernel[3]+tmp[5979]*kernel[4]+tmp[5980]*kernel[5]+tmp[6078]*kernel[6]+tmp[6079]*kernel[7]+tmp[6080]*kernel[8];
				ans[5980]<=tmp[5879]*kernel[0]+tmp[5880]*kernel[1]+tmp[5881]*kernel[2]+tmp[5979]*kernel[3]+tmp[5980]*kernel[4]+tmp[5981]*kernel[5]+tmp[6079]*kernel[6]+tmp[6080]*kernel[7]+tmp[6081]*kernel[8];
				ans[5981]<=tmp[5880]*kernel[0]+tmp[5881]*kernel[1]+tmp[5882]*kernel[2]+tmp[5980]*kernel[3]+tmp[5981]*kernel[4]+tmp[5982]*kernel[5]+tmp[6080]*kernel[6]+tmp[6081]*kernel[7]+tmp[6082]*kernel[8];
				ans[5982]<=tmp[5881]*kernel[0]+tmp[5882]*kernel[1]+tmp[5883]*kernel[2]+tmp[5981]*kernel[3]+tmp[5982]*kernel[4]+tmp[5983]*kernel[5]+tmp[6081]*kernel[6]+tmp[6082]*kernel[7]+tmp[6083]*kernel[8];
				ans[5983]<=tmp[5882]*kernel[0]+tmp[5883]*kernel[1]+tmp[5884]*kernel[2]+tmp[5982]*kernel[3]+tmp[5983]*kernel[4]+tmp[5984]*kernel[5]+tmp[6082]*kernel[6]+tmp[6083]*kernel[7]+tmp[6084]*kernel[8];
				ans[5984]<=tmp[5883]*kernel[0]+tmp[5884]*kernel[1]+tmp[5885]*kernel[2]+tmp[5983]*kernel[3]+tmp[5984]*kernel[4]+tmp[5985]*kernel[5]+tmp[6083]*kernel[6]+tmp[6084]*kernel[7]+tmp[6085]*kernel[8];
				ans[5985]<=tmp[5884]*kernel[0]+tmp[5885]*kernel[1]+tmp[5886]*kernel[2]+tmp[5984]*kernel[3]+tmp[5985]*kernel[4]+tmp[5986]*kernel[5]+tmp[6084]*kernel[6]+tmp[6085]*kernel[7]+tmp[6086]*kernel[8];
				ans[5986]<=tmp[5885]*kernel[0]+tmp[5886]*kernel[1]+tmp[5887]*kernel[2]+tmp[5985]*kernel[3]+tmp[5986]*kernel[4]+tmp[5987]*kernel[5]+tmp[6085]*kernel[6]+tmp[6086]*kernel[7]+tmp[6087]*kernel[8];
				ans[5987]<=tmp[5886]*kernel[0]+tmp[5887]*kernel[1]+tmp[5888]*kernel[2]+tmp[5986]*kernel[3]+tmp[5987]*kernel[4]+tmp[5988]*kernel[5]+tmp[6086]*kernel[6]+tmp[6087]*kernel[7]+tmp[6088]*kernel[8];
				ans[5988]<=tmp[5887]*kernel[0]+tmp[5888]*kernel[1]+tmp[5889]*kernel[2]+tmp[5987]*kernel[3]+tmp[5988]*kernel[4]+tmp[5989]*kernel[5]+tmp[6087]*kernel[6]+tmp[6088]*kernel[7]+tmp[6089]*kernel[8];
				ans[5989]<=tmp[5888]*kernel[0]+tmp[5889]*kernel[1]+tmp[5890]*kernel[2]+tmp[5988]*kernel[3]+tmp[5989]*kernel[4]+tmp[5990]*kernel[5]+tmp[6088]*kernel[6]+tmp[6089]*kernel[7]+tmp[6090]*kernel[8];
				ans[5990]<=tmp[5889]*kernel[0]+tmp[5890]*kernel[1]+tmp[5891]*kernel[2]+tmp[5989]*kernel[3]+tmp[5990]*kernel[4]+tmp[5991]*kernel[5]+tmp[6089]*kernel[6]+tmp[6090]*kernel[7]+tmp[6091]*kernel[8];
				ans[5991]<=tmp[5890]*kernel[0]+tmp[5891]*kernel[1]+tmp[5892]*kernel[2]+tmp[5990]*kernel[3]+tmp[5991]*kernel[4]+tmp[5992]*kernel[5]+tmp[6090]*kernel[6]+tmp[6091]*kernel[7]+tmp[6092]*kernel[8];
				ans[5992]<=tmp[5891]*kernel[0]+tmp[5892]*kernel[1]+tmp[5893]*kernel[2]+tmp[5991]*kernel[3]+tmp[5992]*kernel[4]+tmp[5993]*kernel[5]+tmp[6091]*kernel[6]+tmp[6092]*kernel[7]+tmp[6093]*kernel[8];
				ans[5993]<=tmp[5892]*kernel[0]+tmp[5893]*kernel[1]+tmp[5894]*kernel[2]+tmp[5992]*kernel[3]+tmp[5993]*kernel[4]+tmp[5994]*kernel[5]+tmp[6092]*kernel[6]+tmp[6093]*kernel[7]+tmp[6094]*kernel[8];
				ans[5994]<=tmp[5893]*kernel[0]+tmp[5894]*kernel[1]+tmp[5895]*kernel[2]+tmp[5993]*kernel[3]+tmp[5994]*kernel[4]+tmp[5995]*kernel[5]+tmp[6093]*kernel[6]+tmp[6094]*kernel[7]+tmp[6095]*kernel[8];
				ans[5995]<=tmp[5894]*kernel[0]+tmp[5895]*kernel[1]+tmp[5896]*kernel[2]+tmp[5994]*kernel[3]+tmp[5995]*kernel[4]+tmp[5996]*kernel[5]+tmp[6094]*kernel[6]+tmp[6095]*kernel[7]+tmp[6096]*kernel[8];
				ans[5996]<=tmp[5895]*kernel[0]+tmp[5896]*kernel[1]+tmp[5897]*kernel[2]+tmp[5995]*kernel[3]+tmp[5996]*kernel[4]+tmp[5997]*kernel[5]+tmp[6095]*kernel[6]+tmp[6096]*kernel[7]+tmp[6097]*kernel[8];
				ans[5997]<=tmp[5896]*kernel[0]+tmp[5897]*kernel[1]+tmp[5898]*kernel[2]+tmp[5996]*kernel[3]+tmp[5997]*kernel[4]+tmp[5998]*kernel[5]+tmp[6096]*kernel[6]+tmp[6097]*kernel[7]+tmp[6098]*kernel[8];
				ans[5998]<=tmp[5897]*kernel[0]+tmp[5898]*kernel[1]+tmp[5899]*kernel[2]+tmp[5997]*kernel[3]+tmp[5998]*kernel[4]+tmp[5999]*kernel[5]+tmp[6097]*kernel[6]+tmp[6098]*kernel[7]+tmp[6099]*kernel[8];
				ans[5999]<=tmp[5898]*kernel[0]+tmp[5899]*kernel[1]+tmp[5998]*kernel[3]+tmp[5999]*kernel[4]+tmp[6098]*kernel[6]+tmp[6099]*kernel[7];
				ans[6000]<=tmp[5900]*kernel[1]+tmp[5901]*kernel[2]+tmp[6000]*kernel[4]+tmp[6001]*kernel[5]+tmp[6100]*kernel[7]+tmp[6101]*kernel[8];
				ans[6001]<=tmp[5900]*kernel[0]+tmp[5901]*kernel[1]+tmp[5902]*kernel[2]+tmp[6000]*kernel[3]+tmp[6001]*kernel[4]+tmp[6002]*kernel[5]+tmp[6100]*kernel[6]+tmp[6101]*kernel[7]+tmp[6102]*kernel[8];
				ans[6002]<=tmp[5901]*kernel[0]+tmp[5902]*kernel[1]+tmp[5903]*kernel[2]+tmp[6001]*kernel[3]+tmp[6002]*kernel[4]+tmp[6003]*kernel[5]+tmp[6101]*kernel[6]+tmp[6102]*kernel[7]+tmp[6103]*kernel[8];
				ans[6003]<=tmp[5902]*kernel[0]+tmp[5903]*kernel[1]+tmp[5904]*kernel[2]+tmp[6002]*kernel[3]+tmp[6003]*kernel[4]+tmp[6004]*kernel[5]+tmp[6102]*kernel[6]+tmp[6103]*kernel[7]+tmp[6104]*kernel[8];
				ans[6004]<=tmp[5903]*kernel[0]+tmp[5904]*kernel[1]+tmp[5905]*kernel[2]+tmp[6003]*kernel[3]+tmp[6004]*kernel[4]+tmp[6005]*kernel[5]+tmp[6103]*kernel[6]+tmp[6104]*kernel[7]+tmp[6105]*kernel[8];
				ans[6005]<=tmp[5904]*kernel[0]+tmp[5905]*kernel[1]+tmp[5906]*kernel[2]+tmp[6004]*kernel[3]+tmp[6005]*kernel[4]+tmp[6006]*kernel[5]+tmp[6104]*kernel[6]+tmp[6105]*kernel[7]+tmp[6106]*kernel[8];
				ans[6006]<=tmp[5905]*kernel[0]+tmp[5906]*kernel[1]+tmp[5907]*kernel[2]+tmp[6005]*kernel[3]+tmp[6006]*kernel[4]+tmp[6007]*kernel[5]+tmp[6105]*kernel[6]+tmp[6106]*kernel[7]+tmp[6107]*kernel[8];
				ans[6007]<=tmp[5906]*kernel[0]+tmp[5907]*kernel[1]+tmp[5908]*kernel[2]+tmp[6006]*kernel[3]+tmp[6007]*kernel[4]+tmp[6008]*kernel[5]+tmp[6106]*kernel[6]+tmp[6107]*kernel[7]+tmp[6108]*kernel[8];
				ans[6008]<=tmp[5907]*kernel[0]+tmp[5908]*kernel[1]+tmp[5909]*kernel[2]+tmp[6007]*kernel[3]+tmp[6008]*kernel[4]+tmp[6009]*kernel[5]+tmp[6107]*kernel[6]+tmp[6108]*kernel[7]+tmp[6109]*kernel[8];
				ans[6009]<=tmp[5908]*kernel[0]+tmp[5909]*kernel[1]+tmp[5910]*kernel[2]+tmp[6008]*kernel[3]+tmp[6009]*kernel[4]+tmp[6010]*kernel[5]+tmp[6108]*kernel[6]+tmp[6109]*kernel[7]+tmp[6110]*kernel[8];
				ans[6010]<=tmp[5909]*kernel[0]+tmp[5910]*kernel[1]+tmp[5911]*kernel[2]+tmp[6009]*kernel[3]+tmp[6010]*kernel[4]+tmp[6011]*kernel[5]+tmp[6109]*kernel[6]+tmp[6110]*kernel[7]+tmp[6111]*kernel[8];
				ans[6011]<=tmp[5910]*kernel[0]+tmp[5911]*kernel[1]+tmp[5912]*kernel[2]+tmp[6010]*kernel[3]+tmp[6011]*kernel[4]+tmp[6012]*kernel[5]+tmp[6110]*kernel[6]+tmp[6111]*kernel[7]+tmp[6112]*kernel[8];
				ans[6012]<=tmp[5911]*kernel[0]+tmp[5912]*kernel[1]+tmp[5913]*kernel[2]+tmp[6011]*kernel[3]+tmp[6012]*kernel[4]+tmp[6013]*kernel[5]+tmp[6111]*kernel[6]+tmp[6112]*kernel[7]+tmp[6113]*kernel[8];
				ans[6013]<=tmp[5912]*kernel[0]+tmp[5913]*kernel[1]+tmp[5914]*kernel[2]+tmp[6012]*kernel[3]+tmp[6013]*kernel[4]+tmp[6014]*kernel[5]+tmp[6112]*kernel[6]+tmp[6113]*kernel[7]+tmp[6114]*kernel[8];
				ans[6014]<=tmp[5913]*kernel[0]+tmp[5914]*kernel[1]+tmp[5915]*kernel[2]+tmp[6013]*kernel[3]+tmp[6014]*kernel[4]+tmp[6015]*kernel[5]+tmp[6113]*kernel[6]+tmp[6114]*kernel[7]+tmp[6115]*kernel[8];
				ans[6015]<=tmp[5914]*kernel[0]+tmp[5915]*kernel[1]+tmp[5916]*kernel[2]+tmp[6014]*kernel[3]+tmp[6015]*kernel[4]+tmp[6016]*kernel[5]+tmp[6114]*kernel[6]+tmp[6115]*kernel[7]+tmp[6116]*kernel[8];
				ans[6016]<=tmp[5915]*kernel[0]+tmp[5916]*kernel[1]+tmp[5917]*kernel[2]+tmp[6015]*kernel[3]+tmp[6016]*kernel[4]+tmp[6017]*kernel[5]+tmp[6115]*kernel[6]+tmp[6116]*kernel[7]+tmp[6117]*kernel[8];
				ans[6017]<=tmp[5916]*kernel[0]+tmp[5917]*kernel[1]+tmp[5918]*kernel[2]+tmp[6016]*kernel[3]+tmp[6017]*kernel[4]+tmp[6018]*kernel[5]+tmp[6116]*kernel[6]+tmp[6117]*kernel[7]+tmp[6118]*kernel[8];
				ans[6018]<=tmp[5917]*kernel[0]+tmp[5918]*kernel[1]+tmp[5919]*kernel[2]+tmp[6017]*kernel[3]+tmp[6018]*kernel[4]+tmp[6019]*kernel[5]+tmp[6117]*kernel[6]+tmp[6118]*kernel[7]+tmp[6119]*kernel[8];
				ans[6019]<=tmp[5918]*kernel[0]+tmp[5919]*kernel[1]+tmp[5920]*kernel[2]+tmp[6018]*kernel[3]+tmp[6019]*kernel[4]+tmp[6020]*kernel[5]+tmp[6118]*kernel[6]+tmp[6119]*kernel[7]+tmp[6120]*kernel[8];
				ans[6020]<=tmp[5919]*kernel[0]+tmp[5920]*kernel[1]+tmp[5921]*kernel[2]+tmp[6019]*kernel[3]+tmp[6020]*kernel[4]+tmp[6021]*kernel[5]+tmp[6119]*kernel[6]+tmp[6120]*kernel[7]+tmp[6121]*kernel[8];
				ans[6021]<=tmp[5920]*kernel[0]+tmp[5921]*kernel[1]+tmp[5922]*kernel[2]+tmp[6020]*kernel[3]+tmp[6021]*kernel[4]+tmp[6022]*kernel[5]+tmp[6120]*kernel[6]+tmp[6121]*kernel[7]+tmp[6122]*kernel[8];
				ans[6022]<=tmp[5921]*kernel[0]+tmp[5922]*kernel[1]+tmp[5923]*kernel[2]+tmp[6021]*kernel[3]+tmp[6022]*kernel[4]+tmp[6023]*kernel[5]+tmp[6121]*kernel[6]+tmp[6122]*kernel[7]+tmp[6123]*kernel[8];
				ans[6023]<=tmp[5922]*kernel[0]+tmp[5923]*kernel[1]+tmp[5924]*kernel[2]+tmp[6022]*kernel[3]+tmp[6023]*kernel[4]+tmp[6024]*kernel[5]+tmp[6122]*kernel[6]+tmp[6123]*kernel[7]+tmp[6124]*kernel[8];
				ans[6024]<=tmp[5923]*kernel[0]+tmp[5924]*kernel[1]+tmp[5925]*kernel[2]+tmp[6023]*kernel[3]+tmp[6024]*kernel[4]+tmp[6025]*kernel[5]+tmp[6123]*kernel[6]+tmp[6124]*kernel[7]+tmp[6125]*kernel[8];
				ans[6025]<=tmp[5924]*kernel[0]+tmp[5925]*kernel[1]+tmp[5926]*kernel[2]+tmp[6024]*kernel[3]+tmp[6025]*kernel[4]+tmp[6026]*kernel[5]+tmp[6124]*kernel[6]+tmp[6125]*kernel[7]+tmp[6126]*kernel[8];
				ans[6026]<=tmp[5925]*kernel[0]+tmp[5926]*kernel[1]+tmp[5927]*kernel[2]+tmp[6025]*kernel[3]+tmp[6026]*kernel[4]+tmp[6027]*kernel[5]+tmp[6125]*kernel[6]+tmp[6126]*kernel[7]+tmp[6127]*kernel[8];
				ans[6027]<=tmp[5926]*kernel[0]+tmp[5927]*kernel[1]+tmp[5928]*kernel[2]+tmp[6026]*kernel[3]+tmp[6027]*kernel[4]+tmp[6028]*kernel[5]+tmp[6126]*kernel[6]+tmp[6127]*kernel[7]+tmp[6128]*kernel[8];
				ans[6028]<=tmp[5927]*kernel[0]+tmp[5928]*kernel[1]+tmp[5929]*kernel[2]+tmp[6027]*kernel[3]+tmp[6028]*kernel[4]+tmp[6029]*kernel[5]+tmp[6127]*kernel[6]+tmp[6128]*kernel[7]+tmp[6129]*kernel[8];
				ans[6029]<=tmp[5928]*kernel[0]+tmp[5929]*kernel[1]+tmp[5930]*kernel[2]+tmp[6028]*kernel[3]+tmp[6029]*kernel[4]+tmp[6030]*kernel[5]+tmp[6128]*kernel[6]+tmp[6129]*kernel[7]+tmp[6130]*kernel[8];
				ans[6030]<=tmp[5929]*kernel[0]+tmp[5930]*kernel[1]+tmp[5931]*kernel[2]+tmp[6029]*kernel[3]+tmp[6030]*kernel[4]+tmp[6031]*kernel[5]+tmp[6129]*kernel[6]+tmp[6130]*kernel[7]+tmp[6131]*kernel[8];
				ans[6031]<=tmp[5930]*kernel[0]+tmp[5931]*kernel[1]+tmp[5932]*kernel[2]+tmp[6030]*kernel[3]+tmp[6031]*kernel[4]+tmp[6032]*kernel[5]+tmp[6130]*kernel[6]+tmp[6131]*kernel[7]+tmp[6132]*kernel[8];
				ans[6032]<=tmp[5931]*kernel[0]+tmp[5932]*kernel[1]+tmp[5933]*kernel[2]+tmp[6031]*kernel[3]+tmp[6032]*kernel[4]+tmp[6033]*kernel[5]+tmp[6131]*kernel[6]+tmp[6132]*kernel[7]+tmp[6133]*kernel[8];
				ans[6033]<=tmp[5932]*kernel[0]+tmp[5933]*kernel[1]+tmp[5934]*kernel[2]+tmp[6032]*kernel[3]+tmp[6033]*kernel[4]+tmp[6034]*kernel[5]+tmp[6132]*kernel[6]+tmp[6133]*kernel[7]+tmp[6134]*kernel[8];
				ans[6034]<=tmp[5933]*kernel[0]+tmp[5934]*kernel[1]+tmp[5935]*kernel[2]+tmp[6033]*kernel[3]+tmp[6034]*kernel[4]+tmp[6035]*kernel[5]+tmp[6133]*kernel[6]+tmp[6134]*kernel[7]+tmp[6135]*kernel[8];
				ans[6035]<=tmp[5934]*kernel[0]+tmp[5935]*kernel[1]+tmp[5936]*kernel[2]+tmp[6034]*kernel[3]+tmp[6035]*kernel[4]+tmp[6036]*kernel[5]+tmp[6134]*kernel[6]+tmp[6135]*kernel[7]+tmp[6136]*kernel[8];
				ans[6036]<=tmp[5935]*kernel[0]+tmp[5936]*kernel[1]+tmp[5937]*kernel[2]+tmp[6035]*kernel[3]+tmp[6036]*kernel[4]+tmp[6037]*kernel[5]+tmp[6135]*kernel[6]+tmp[6136]*kernel[7]+tmp[6137]*kernel[8];
				ans[6037]<=tmp[5936]*kernel[0]+tmp[5937]*kernel[1]+tmp[5938]*kernel[2]+tmp[6036]*kernel[3]+tmp[6037]*kernel[4]+tmp[6038]*kernel[5]+tmp[6136]*kernel[6]+tmp[6137]*kernel[7]+tmp[6138]*kernel[8];
				ans[6038]<=tmp[5937]*kernel[0]+tmp[5938]*kernel[1]+tmp[5939]*kernel[2]+tmp[6037]*kernel[3]+tmp[6038]*kernel[4]+tmp[6039]*kernel[5]+tmp[6137]*kernel[6]+tmp[6138]*kernel[7]+tmp[6139]*kernel[8];
				ans[6039]<=tmp[5938]*kernel[0]+tmp[5939]*kernel[1]+tmp[5940]*kernel[2]+tmp[6038]*kernel[3]+tmp[6039]*kernel[4]+tmp[6040]*kernel[5]+tmp[6138]*kernel[6]+tmp[6139]*kernel[7]+tmp[6140]*kernel[8];
				ans[6040]<=tmp[5939]*kernel[0]+tmp[5940]*kernel[1]+tmp[5941]*kernel[2]+tmp[6039]*kernel[3]+tmp[6040]*kernel[4]+tmp[6041]*kernel[5]+tmp[6139]*kernel[6]+tmp[6140]*kernel[7]+tmp[6141]*kernel[8];
				ans[6041]<=tmp[5940]*kernel[0]+tmp[5941]*kernel[1]+tmp[5942]*kernel[2]+tmp[6040]*kernel[3]+tmp[6041]*kernel[4]+tmp[6042]*kernel[5]+tmp[6140]*kernel[6]+tmp[6141]*kernel[7]+tmp[6142]*kernel[8];
				ans[6042]<=tmp[5941]*kernel[0]+tmp[5942]*kernel[1]+tmp[5943]*kernel[2]+tmp[6041]*kernel[3]+tmp[6042]*kernel[4]+tmp[6043]*kernel[5]+tmp[6141]*kernel[6]+tmp[6142]*kernel[7]+tmp[6143]*kernel[8];
				ans[6043]<=tmp[5942]*kernel[0]+tmp[5943]*kernel[1]+tmp[5944]*kernel[2]+tmp[6042]*kernel[3]+tmp[6043]*kernel[4]+tmp[6044]*kernel[5]+tmp[6142]*kernel[6]+tmp[6143]*kernel[7]+tmp[6144]*kernel[8];
				ans[6044]<=tmp[5943]*kernel[0]+tmp[5944]*kernel[1]+tmp[5945]*kernel[2]+tmp[6043]*kernel[3]+tmp[6044]*kernel[4]+tmp[6045]*kernel[5]+tmp[6143]*kernel[6]+tmp[6144]*kernel[7]+tmp[6145]*kernel[8];
				ans[6045]<=tmp[5944]*kernel[0]+tmp[5945]*kernel[1]+tmp[5946]*kernel[2]+tmp[6044]*kernel[3]+tmp[6045]*kernel[4]+tmp[6046]*kernel[5]+tmp[6144]*kernel[6]+tmp[6145]*kernel[7]+tmp[6146]*kernel[8];
				ans[6046]<=tmp[5945]*kernel[0]+tmp[5946]*kernel[1]+tmp[5947]*kernel[2]+tmp[6045]*kernel[3]+tmp[6046]*kernel[4]+tmp[6047]*kernel[5]+tmp[6145]*kernel[6]+tmp[6146]*kernel[7]+tmp[6147]*kernel[8];
				ans[6047]<=tmp[5946]*kernel[0]+tmp[5947]*kernel[1]+tmp[5948]*kernel[2]+tmp[6046]*kernel[3]+tmp[6047]*kernel[4]+tmp[6048]*kernel[5]+tmp[6146]*kernel[6]+tmp[6147]*kernel[7]+tmp[6148]*kernel[8];
				ans[6048]<=tmp[5947]*kernel[0]+tmp[5948]*kernel[1]+tmp[5949]*kernel[2]+tmp[6047]*kernel[3]+tmp[6048]*kernel[4]+tmp[6049]*kernel[5]+tmp[6147]*kernel[6]+tmp[6148]*kernel[7]+tmp[6149]*kernel[8];
				ans[6049]<=tmp[5948]*kernel[0]+tmp[5949]*kernel[1]+tmp[5950]*kernel[2]+tmp[6048]*kernel[3]+tmp[6049]*kernel[4]+tmp[6050]*kernel[5]+tmp[6148]*kernel[6]+tmp[6149]*kernel[7]+tmp[6150]*kernel[8];
				ans[6050]<=tmp[5949]*kernel[0]+tmp[5950]*kernel[1]+tmp[5951]*kernel[2]+tmp[6049]*kernel[3]+tmp[6050]*kernel[4]+tmp[6051]*kernel[5]+tmp[6149]*kernel[6]+tmp[6150]*kernel[7]+tmp[6151]*kernel[8];
				ans[6051]<=tmp[5950]*kernel[0]+tmp[5951]*kernel[1]+tmp[5952]*kernel[2]+tmp[6050]*kernel[3]+tmp[6051]*kernel[4]+tmp[6052]*kernel[5]+tmp[6150]*kernel[6]+tmp[6151]*kernel[7]+tmp[6152]*kernel[8];
				ans[6052]<=tmp[5951]*kernel[0]+tmp[5952]*kernel[1]+tmp[5953]*kernel[2]+tmp[6051]*kernel[3]+tmp[6052]*kernel[4]+tmp[6053]*kernel[5]+tmp[6151]*kernel[6]+tmp[6152]*kernel[7]+tmp[6153]*kernel[8];
				ans[6053]<=tmp[5952]*kernel[0]+tmp[5953]*kernel[1]+tmp[5954]*kernel[2]+tmp[6052]*kernel[3]+tmp[6053]*kernel[4]+tmp[6054]*kernel[5]+tmp[6152]*kernel[6]+tmp[6153]*kernel[7]+tmp[6154]*kernel[8];
				ans[6054]<=tmp[5953]*kernel[0]+tmp[5954]*kernel[1]+tmp[5955]*kernel[2]+tmp[6053]*kernel[3]+tmp[6054]*kernel[4]+tmp[6055]*kernel[5]+tmp[6153]*kernel[6]+tmp[6154]*kernel[7]+tmp[6155]*kernel[8];
				ans[6055]<=tmp[5954]*kernel[0]+tmp[5955]*kernel[1]+tmp[5956]*kernel[2]+tmp[6054]*kernel[3]+tmp[6055]*kernel[4]+tmp[6056]*kernel[5]+tmp[6154]*kernel[6]+tmp[6155]*kernel[7]+tmp[6156]*kernel[8];
				ans[6056]<=tmp[5955]*kernel[0]+tmp[5956]*kernel[1]+tmp[5957]*kernel[2]+tmp[6055]*kernel[3]+tmp[6056]*kernel[4]+tmp[6057]*kernel[5]+tmp[6155]*kernel[6]+tmp[6156]*kernel[7]+tmp[6157]*kernel[8];
				ans[6057]<=tmp[5956]*kernel[0]+tmp[5957]*kernel[1]+tmp[5958]*kernel[2]+tmp[6056]*kernel[3]+tmp[6057]*kernel[4]+tmp[6058]*kernel[5]+tmp[6156]*kernel[6]+tmp[6157]*kernel[7]+tmp[6158]*kernel[8];
				ans[6058]<=tmp[5957]*kernel[0]+tmp[5958]*kernel[1]+tmp[5959]*kernel[2]+tmp[6057]*kernel[3]+tmp[6058]*kernel[4]+tmp[6059]*kernel[5]+tmp[6157]*kernel[6]+tmp[6158]*kernel[7]+tmp[6159]*kernel[8];
				ans[6059]<=tmp[5958]*kernel[0]+tmp[5959]*kernel[1]+tmp[5960]*kernel[2]+tmp[6058]*kernel[3]+tmp[6059]*kernel[4]+tmp[6060]*kernel[5]+tmp[6158]*kernel[6]+tmp[6159]*kernel[7]+tmp[6160]*kernel[8];
				ans[6060]<=tmp[5959]*kernel[0]+tmp[5960]*kernel[1]+tmp[5961]*kernel[2]+tmp[6059]*kernel[3]+tmp[6060]*kernel[4]+tmp[6061]*kernel[5]+tmp[6159]*kernel[6]+tmp[6160]*kernel[7]+tmp[6161]*kernel[8];
				ans[6061]<=tmp[5960]*kernel[0]+tmp[5961]*kernel[1]+tmp[5962]*kernel[2]+tmp[6060]*kernel[3]+tmp[6061]*kernel[4]+tmp[6062]*kernel[5]+tmp[6160]*kernel[6]+tmp[6161]*kernel[7]+tmp[6162]*kernel[8];
				ans[6062]<=tmp[5961]*kernel[0]+tmp[5962]*kernel[1]+tmp[5963]*kernel[2]+tmp[6061]*kernel[3]+tmp[6062]*kernel[4]+tmp[6063]*kernel[5]+tmp[6161]*kernel[6]+tmp[6162]*kernel[7]+tmp[6163]*kernel[8];
				ans[6063]<=tmp[5962]*kernel[0]+tmp[5963]*kernel[1]+tmp[5964]*kernel[2]+tmp[6062]*kernel[3]+tmp[6063]*kernel[4]+tmp[6064]*kernel[5]+tmp[6162]*kernel[6]+tmp[6163]*kernel[7]+tmp[6164]*kernel[8];
				ans[6064]<=tmp[5963]*kernel[0]+tmp[5964]*kernel[1]+tmp[5965]*kernel[2]+tmp[6063]*kernel[3]+tmp[6064]*kernel[4]+tmp[6065]*kernel[5]+tmp[6163]*kernel[6]+tmp[6164]*kernel[7]+tmp[6165]*kernel[8];
				ans[6065]<=tmp[5964]*kernel[0]+tmp[5965]*kernel[1]+tmp[5966]*kernel[2]+tmp[6064]*kernel[3]+tmp[6065]*kernel[4]+tmp[6066]*kernel[5]+tmp[6164]*kernel[6]+tmp[6165]*kernel[7]+tmp[6166]*kernel[8];
				ans[6066]<=tmp[5965]*kernel[0]+tmp[5966]*kernel[1]+tmp[5967]*kernel[2]+tmp[6065]*kernel[3]+tmp[6066]*kernel[4]+tmp[6067]*kernel[5]+tmp[6165]*kernel[6]+tmp[6166]*kernel[7]+tmp[6167]*kernel[8];
				ans[6067]<=tmp[5966]*kernel[0]+tmp[5967]*kernel[1]+tmp[5968]*kernel[2]+tmp[6066]*kernel[3]+tmp[6067]*kernel[4]+tmp[6068]*kernel[5]+tmp[6166]*kernel[6]+tmp[6167]*kernel[7]+tmp[6168]*kernel[8];
				ans[6068]<=tmp[5967]*kernel[0]+tmp[5968]*kernel[1]+tmp[5969]*kernel[2]+tmp[6067]*kernel[3]+tmp[6068]*kernel[4]+tmp[6069]*kernel[5]+tmp[6167]*kernel[6]+tmp[6168]*kernel[7]+tmp[6169]*kernel[8];
				ans[6069]<=tmp[5968]*kernel[0]+tmp[5969]*kernel[1]+tmp[5970]*kernel[2]+tmp[6068]*kernel[3]+tmp[6069]*kernel[4]+tmp[6070]*kernel[5]+tmp[6168]*kernel[6]+tmp[6169]*kernel[7]+tmp[6170]*kernel[8];
				ans[6070]<=tmp[5969]*kernel[0]+tmp[5970]*kernel[1]+tmp[5971]*kernel[2]+tmp[6069]*kernel[3]+tmp[6070]*kernel[4]+tmp[6071]*kernel[5]+tmp[6169]*kernel[6]+tmp[6170]*kernel[7]+tmp[6171]*kernel[8];
				ans[6071]<=tmp[5970]*kernel[0]+tmp[5971]*kernel[1]+tmp[5972]*kernel[2]+tmp[6070]*kernel[3]+tmp[6071]*kernel[4]+tmp[6072]*kernel[5]+tmp[6170]*kernel[6]+tmp[6171]*kernel[7]+tmp[6172]*kernel[8];
				ans[6072]<=tmp[5971]*kernel[0]+tmp[5972]*kernel[1]+tmp[5973]*kernel[2]+tmp[6071]*kernel[3]+tmp[6072]*kernel[4]+tmp[6073]*kernel[5]+tmp[6171]*kernel[6]+tmp[6172]*kernel[7]+tmp[6173]*kernel[8];
				ans[6073]<=tmp[5972]*kernel[0]+tmp[5973]*kernel[1]+tmp[5974]*kernel[2]+tmp[6072]*kernel[3]+tmp[6073]*kernel[4]+tmp[6074]*kernel[5]+tmp[6172]*kernel[6]+tmp[6173]*kernel[7]+tmp[6174]*kernel[8];
				ans[6074]<=tmp[5973]*kernel[0]+tmp[5974]*kernel[1]+tmp[5975]*kernel[2]+tmp[6073]*kernel[3]+tmp[6074]*kernel[4]+tmp[6075]*kernel[5]+tmp[6173]*kernel[6]+tmp[6174]*kernel[7]+tmp[6175]*kernel[8];
				ans[6075]<=tmp[5974]*kernel[0]+tmp[5975]*kernel[1]+tmp[5976]*kernel[2]+tmp[6074]*kernel[3]+tmp[6075]*kernel[4]+tmp[6076]*kernel[5]+tmp[6174]*kernel[6]+tmp[6175]*kernel[7]+tmp[6176]*kernel[8];
				ans[6076]<=tmp[5975]*kernel[0]+tmp[5976]*kernel[1]+tmp[5977]*kernel[2]+tmp[6075]*kernel[3]+tmp[6076]*kernel[4]+tmp[6077]*kernel[5]+tmp[6175]*kernel[6]+tmp[6176]*kernel[7]+tmp[6177]*kernel[8];
				ans[6077]<=tmp[5976]*kernel[0]+tmp[5977]*kernel[1]+tmp[5978]*kernel[2]+tmp[6076]*kernel[3]+tmp[6077]*kernel[4]+tmp[6078]*kernel[5]+tmp[6176]*kernel[6]+tmp[6177]*kernel[7]+tmp[6178]*kernel[8];
				ans[6078]<=tmp[5977]*kernel[0]+tmp[5978]*kernel[1]+tmp[5979]*kernel[2]+tmp[6077]*kernel[3]+tmp[6078]*kernel[4]+tmp[6079]*kernel[5]+tmp[6177]*kernel[6]+tmp[6178]*kernel[7]+tmp[6179]*kernel[8];
				ans[6079]<=tmp[5978]*kernel[0]+tmp[5979]*kernel[1]+tmp[5980]*kernel[2]+tmp[6078]*kernel[3]+tmp[6079]*kernel[4]+tmp[6080]*kernel[5]+tmp[6178]*kernel[6]+tmp[6179]*kernel[7]+tmp[6180]*kernel[8];
				ans[6080]<=tmp[5979]*kernel[0]+tmp[5980]*kernel[1]+tmp[5981]*kernel[2]+tmp[6079]*kernel[3]+tmp[6080]*kernel[4]+tmp[6081]*kernel[5]+tmp[6179]*kernel[6]+tmp[6180]*kernel[7]+tmp[6181]*kernel[8];
				ans[6081]<=tmp[5980]*kernel[0]+tmp[5981]*kernel[1]+tmp[5982]*kernel[2]+tmp[6080]*kernel[3]+tmp[6081]*kernel[4]+tmp[6082]*kernel[5]+tmp[6180]*kernel[6]+tmp[6181]*kernel[7]+tmp[6182]*kernel[8];
				ans[6082]<=tmp[5981]*kernel[0]+tmp[5982]*kernel[1]+tmp[5983]*kernel[2]+tmp[6081]*kernel[3]+tmp[6082]*kernel[4]+tmp[6083]*kernel[5]+tmp[6181]*kernel[6]+tmp[6182]*kernel[7]+tmp[6183]*kernel[8];
				ans[6083]<=tmp[5982]*kernel[0]+tmp[5983]*kernel[1]+tmp[5984]*kernel[2]+tmp[6082]*kernel[3]+tmp[6083]*kernel[4]+tmp[6084]*kernel[5]+tmp[6182]*kernel[6]+tmp[6183]*kernel[7]+tmp[6184]*kernel[8];
				ans[6084]<=tmp[5983]*kernel[0]+tmp[5984]*kernel[1]+tmp[5985]*kernel[2]+tmp[6083]*kernel[3]+tmp[6084]*kernel[4]+tmp[6085]*kernel[5]+tmp[6183]*kernel[6]+tmp[6184]*kernel[7]+tmp[6185]*kernel[8];
				ans[6085]<=tmp[5984]*kernel[0]+tmp[5985]*kernel[1]+tmp[5986]*kernel[2]+tmp[6084]*kernel[3]+tmp[6085]*kernel[4]+tmp[6086]*kernel[5]+tmp[6184]*kernel[6]+tmp[6185]*kernel[7]+tmp[6186]*kernel[8];
				ans[6086]<=tmp[5985]*kernel[0]+tmp[5986]*kernel[1]+tmp[5987]*kernel[2]+tmp[6085]*kernel[3]+tmp[6086]*kernel[4]+tmp[6087]*kernel[5]+tmp[6185]*kernel[6]+tmp[6186]*kernel[7]+tmp[6187]*kernel[8];
				ans[6087]<=tmp[5986]*kernel[0]+tmp[5987]*kernel[1]+tmp[5988]*kernel[2]+tmp[6086]*kernel[3]+tmp[6087]*kernel[4]+tmp[6088]*kernel[5]+tmp[6186]*kernel[6]+tmp[6187]*kernel[7]+tmp[6188]*kernel[8];
				ans[6088]<=tmp[5987]*kernel[0]+tmp[5988]*kernel[1]+tmp[5989]*kernel[2]+tmp[6087]*kernel[3]+tmp[6088]*kernel[4]+tmp[6089]*kernel[5]+tmp[6187]*kernel[6]+tmp[6188]*kernel[7]+tmp[6189]*kernel[8];
				ans[6089]<=tmp[5988]*kernel[0]+tmp[5989]*kernel[1]+tmp[5990]*kernel[2]+tmp[6088]*kernel[3]+tmp[6089]*kernel[4]+tmp[6090]*kernel[5]+tmp[6188]*kernel[6]+tmp[6189]*kernel[7]+tmp[6190]*kernel[8];
				ans[6090]<=tmp[5989]*kernel[0]+tmp[5990]*kernel[1]+tmp[5991]*kernel[2]+tmp[6089]*kernel[3]+tmp[6090]*kernel[4]+tmp[6091]*kernel[5]+tmp[6189]*kernel[6]+tmp[6190]*kernel[7]+tmp[6191]*kernel[8];
				ans[6091]<=tmp[5990]*kernel[0]+tmp[5991]*kernel[1]+tmp[5992]*kernel[2]+tmp[6090]*kernel[3]+tmp[6091]*kernel[4]+tmp[6092]*kernel[5]+tmp[6190]*kernel[6]+tmp[6191]*kernel[7]+tmp[6192]*kernel[8];
				ans[6092]<=tmp[5991]*kernel[0]+tmp[5992]*kernel[1]+tmp[5993]*kernel[2]+tmp[6091]*kernel[3]+tmp[6092]*kernel[4]+tmp[6093]*kernel[5]+tmp[6191]*kernel[6]+tmp[6192]*kernel[7]+tmp[6193]*kernel[8];
				ans[6093]<=tmp[5992]*kernel[0]+tmp[5993]*kernel[1]+tmp[5994]*kernel[2]+tmp[6092]*kernel[3]+tmp[6093]*kernel[4]+tmp[6094]*kernel[5]+tmp[6192]*kernel[6]+tmp[6193]*kernel[7]+tmp[6194]*kernel[8];
				ans[6094]<=tmp[5993]*kernel[0]+tmp[5994]*kernel[1]+tmp[5995]*kernel[2]+tmp[6093]*kernel[3]+tmp[6094]*kernel[4]+tmp[6095]*kernel[5]+tmp[6193]*kernel[6]+tmp[6194]*kernel[7]+tmp[6195]*kernel[8];
				ans[6095]<=tmp[5994]*kernel[0]+tmp[5995]*kernel[1]+tmp[5996]*kernel[2]+tmp[6094]*kernel[3]+tmp[6095]*kernel[4]+tmp[6096]*kernel[5]+tmp[6194]*kernel[6]+tmp[6195]*kernel[7]+tmp[6196]*kernel[8];
				ans[6096]<=tmp[5995]*kernel[0]+tmp[5996]*kernel[1]+tmp[5997]*kernel[2]+tmp[6095]*kernel[3]+tmp[6096]*kernel[4]+tmp[6097]*kernel[5]+tmp[6195]*kernel[6]+tmp[6196]*kernel[7]+tmp[6197]*kernel[8];
				ans[6097]<=tmp[5996]*kernel[0]+tmp[5997]*kernel[1]+tmp[5998]*kernel[2]+tmp[6096]*kernel[3]+tmp[6097]*kernel[4]+tmp[6098]*kernel[5]+tmp[6196]*kernel[6]+tmp[6197]*kernel[7]+tmp[6198]*kernel[8];
				ans[6098]<=tmp[5997]*kernel[0]+tmp[5998]*kernel[1]+tmp[5999]*kernel[2]+tmp[6097]*kernel[3]+tmp[6098]*kernel[4]+tmp[6099]*kernel[5]+tmp[6197]*kernel[6]+tmp[6198]*kernel[7]+tmp[6199]*kernel[8];
				ans[6099]<=tmp[5998]*kernel[0]+tmp[5999]*kernel[1]+tmp[6098]*kernel[3]+tmp[6099]*kernel[4]+tmp[6198]*kernel[6]+tmp[6199]*kernel[7];
				ans[6100]<=tmp[6000]*kernel[1]+tmp[6001]*kernel[2]+tmp[6100]*kernel[4]+tmp[6101]*kernel[5]+tmp[6200]*kernel[7]+tmp[6201]*kernel[8];
				ans[6101]<=tmp[6000]*kernel[0]+tmp[6001]*kernel[1]+tmp[6002]*kernel[2]+tmp[6100]*kernel[3]+tmp[6101]*kernel[4]+tmp[6102]*kernel[5]+tmp[6200]*kernel[6]+tmp[6201]*kernel[7]+tmp[6202]*kernel[8];
				ans[6102]<=tmp[6001]*kernel[0]+tmp[6002]*kernel[1]+tmp[6003]*kernel[2]+tmp[6101]*kernel[3]+tmp[6102]*kernel[4]+tmp[6103]*kernel[5]+tmp[6201]*kernel[6]+tmp[6202]*kernel[7]+tmp[6203]*kernel[8];
				ans[6103]<=tmp[6002]*kernel[0]+tmp[6003]*kernel[1]+tmp[6004]*kernel[2]+tmp[6102]*kernel[3]+tmp[6103]*kernel[4]+tmp[6104]*kernel[5]+tmp[6202]*kernel[6]+tmp[6203]*kernel[7]+tmp[6204]*kernel[8];
				ans[6104]<=tmp[6003]*kernel[0]+tmp[6004]*kernel[1]+tmp[6005]*kernel[2]+tmp[6103]*kernel[3]+tmp[6104]*kernel[4]+tmp[6105]*kernel[5]+tmp[6203]*kernel[6]+tmp[6204]*kernel[7]+tmp[6205]*kernel[8];
				ans[6105]<=tmp[6004]*kernel[0]+tmp[6005]*kernel[1]+tmp[6006]*kernel[2]+tmp[6104]*kernel[3]+tmp[6105]*kernel[4]+tmp[6106]*kernel[5]+tmp[6204]*kernel[6]+tmp[6205]*kernel[7]+tmp[6206]*kernel[8];
				ans[6106]<=tmp[6005]*kernel[0]+tmp[6006]*kernel[1]+tmp[6007]*kernel[2]+tmp[6105]*kernel[3]+tmp[6106]*kernel[4]+tmp[6107]*kernel[5]+tmp[6205]*kernel[6]+tmp[6206]*kernel[7]+tmp[6207]*kernel[8];
				ans[6107]<=tmp[6006]*kernel[0]+tmp[6007]*kernel[1]+tmp[6008]*kernel[2]+tmp[6106]*kernel[3]+tmp[6107]*kernel[4]+tmp[6108]*kernel[5]+tmp[6206]*kernel[6]+tmp[6207]*kernel[7]+tmp[6208]*kernel[8];
				ans[6108]<=tmp[6007]*kernel[0]+tmp[6008]*kernel[1]+tmp[6009]*kernel[2]+tmp[6107]*kernel[3]+tmp[6108]*kernel[4]+tmp[6109]*kernel[5]+tmp[6207]*kernel[6]+tmp[6208]*kernel[7]+tmp[6209]*kernel[8];
				ans[6109]<=tmp[6008]*kernel[0]+tmp[6009]*kernel[1]+tmp[6010]*kernel[2]+tmp[6108]*kernel[3]+tmp[6109]*kernel[4]+tmp[6110]*kernel[5]+tmp[6208]*kernel[6]+tmp[6209]*kernel[7]+tmp[6210]*kernel[8];
				ans[6110]<=tmp[6009]*kernel[0]+tmp[6010]*kernel[1]+tmp[6011]*kernel[2]+tmp[6109]*kernel[3]+tmp[6110]*kernel[4]+tmp[6111]*kernel[5]+tmp[6209]*kernel[6]+tmp[6210]*kernel[7]+tmp[6211]*kernel[8];
				ans[6111]<=tmp[6010]*kernel[0]+tmp[6011]*kernel[1]+tmp[6012]*kernel[2]+tmp[6110]*kernel[3]+tmp[6111]*kernel[4]+tmp[6112]*kernel[5]+tmp[6210]*kernel[6]+tmp[6211]*kernel[7]+tmp[6212]*kernel[8];
				ans[6112]<=tmp[6011]*kernel[0]+tmp[6012]*kernel[1]+tmp[6013]*kernel[2]+tmp[6111]*kernel[3]+tmp[6112]*kernel[4]+tmp[6113]*kernel[5]+tmp[6211]*kernel[6]+tmp[6212]*kernel[7]+tmp[6213]*kernel[8];
				ans[6113]<=tmp[6012]*kernel[0]+tmp[6013]*kernel[1]+tmp[6014]*kernel[2]+tmp[6112]*kernel[3]+tmp[6113]*kernel[4]+tmp[6114]*kernel[5]+tmp[6212]*kernel[6]+tmp[6213]*kernel[7]+tmp[6214]*kernel[8];
				ans[6114]<=tmp[6013]*kernel[0]+tmp[6014]*kernel[1]+tmp[6015]*kernel[2]+tmp[6113]*kernel[3]+tmp[6114]*kernel[4]+tmp[6115]*kernel[5]+tmp[6213]*kernel[6]+tmp[6214]*kernel[7]+tmp[6215]*kernel[8];
				ans[6115]<=tmp[6014]*kernel[0]+tmp[6015]*kernel[1]+tmp[6016]*kernel[2]+tmp[6114]*kernel[3]+tmp[6115]*kernel[4]+tmp[6116]*kernel[5]+tmp[6214]*kernel[6]+tmp[6215]*kernel[7]+tmp[6216]*kernel[8];
				ans[6116]<=tmp[6015]*kernel[0]+tmp[6016]*kernel[1]+tmp[6017]*kernel[2]+tmp[6115]*kernel[3]+tmp[6116]*kernel[4]+tmp[6117]*kernel[5]+tmp[6215]*kernel[6]+tmp[6216]*kernel[7]+tmp[6217]*kernel[8];
				ans[6117]<=tmp[6016]*kernel[0]+tmp[6017]*kernel[1]+tmp[6018]*kernel[2]+tmp[6116]*kernel[3]+tmp[6117]*kernel[4]+tmp[6118]*kernel[5]+tmp[6216]*kernel[6]+tmp[6217]*kernel[7]+tmp[6218]*kernel[8];
				ans[6118]<=tmp[6017]*kernel[0]+tmp[6018]*kernel[1]+tmp[6019]*kernel[2]+tmp[6117]*kernel[3]+tmp[6118]*kernel[4]+tmp[6119]*kernel[5]+tmp[6217]*kernel[6]+tmp[6218]*kernel[7]+tmp[6219]*kernel[8];
				ans[6119]<=tmp[6018]*kernel[0]+tmp[6019]*kernel[1]+tmp[6020]*kernel[2]+tmp[6118]*kernel[3]+tmp[6119]*kernel[4]+tmp[6120]*kernel[5]+tmp[6218]*kernel[6]+tmp[6219]*kernel[7]+tmp[6220]*kernel[8];
				ans[6120]<=tmp[6019]*kernel[0]+tmp[6020]*kernel[1]+tmp[6021]*kernel[2]+tmp[6119]*kernel[3]+tmp[6120]*kernel[4]+tmp[6121]*kernel[5]+tmp[6219]*kernel[6]+tmp[6220]*kernel[7]+tmp[6221]*kernel[8];
				ans[6121]<=tmp[6020]*kernel[0]+tmp[6021]*kernel[1]+tmp[6022]*kernel[2]+tmp[6120]*kernel[3]+tmp[6121]*kernel[4]+tmp[6122]*kernel[5]+tmp[6220]*kernel[6]+tmp[6221]*kernel[7]+tmp[6222]*kernel[8];
				ans[6122]<=tmp[6021]*kernel[0]+tmp[6022]*kernel[1]+tmp[6023]*kernel[2]+tmp[6121]*kernel[3]+tmp[6122]*kernel[4]+tmp[6123]*kernel[5]+tmp[6221]*kernel[6]+tmp[6222]*kernel[7]+tmp[6223]*kernel[8];
				ans[6123]<=tmp[6022]*kernel[0]+tmp[6023]*kernel[1]+tmp[6024]*kernel[2]+tmp[6122]*kernel[3]+tmp[6123]*kernel[4]+tmp[6124]*kernel[5]+tmp[6222]*kernel[6]+tmp[6223]*kernel[7]+tmp[6224]*kernel[8];
				ans[6124]<=tmp[6023]*kernel[0]+tmp[6024]*kernel[1]+tmp[6025]*kernel[2]+tmp[6123]*kernel[3]+tmp[6124]*kernel[4]+tmp[6125]*kernel[5]+tmp[6223]*kernel[6]+tmp[6224]*kernel[7]+tmp[6225]*kernel[8];
				ans[6125]<=tmp[6024]*kernel[0]+tmp[6025]*kernel[1]+tmp[6026]*kernel[2]+tmp[6124]*kernel[3]+tmp[6125]*kernel[4]+tmp[6126]*kernel[5]+tmp[6224]*kernel[6]+tmp[6225]*kernel[7]+tmp[6226]*kernel[8];
				ans[6126]<=tmp[6025]*kernel[0]+tmp[6026]*kernel[1]+tmp[6027]*kernel[2]+tmp[6125]*kernel[3]+tmp[6126]*kernel[4]+tmp[6127]*kernel[5]+tmp[6225]*kernel[6]+tmp[6226]*kernel[7]+tmp[6227]*kernel[8];
				ans[6127]<=tmp[6026]*kernel[0]+tmp[6027]*kernel[1]+tmp[6028]*kernel[2]+tmp[6126]*kernel[3]+tmp[6127]*kernel[4]+tmp[6128]*kernel[5]+tmp[6226]*kernel[6]+tmp[6227]*kernel[7]+tmp[6228]*kernel[8];
				ans[6128]<=tmp[6027]*kernel[0]+tmp[6028]*kernel[1]+tmp[6029]*kernel[2]+tmp[6127]*kernel[3]+tmp[6128]*kernel[4]+tmp[6129]*kernel[5]+tmp[6227]*kernel[6]+tmp[6228]*kernel[7]+tmp[6229]*kernel[8];
				ans[6129]<=tmp[6028]*kernel[0]+tmp[6029]*kernel[1]+tmp[6030]*kernel[2]+tmp[6128]*kernel[3]+tmp[6129]*kernel[4]+tmp[6130]*kernel[5]+tmp[6228]*kernel[6]+tmp[6229]*kernel[7]+tmp[6230]*kernel[8];
				ans[6130]<=tmp[6029]*kernel[0]+tmp[6030]*kernel[1]+tmp[6031]*kernel[2]+tmp[6129]*kernel[3]+tmp[6130]*kernel[4]+tmp[6131]*kernel[5]+tmp[6229]*kernel[6]+tmp[6230]*kernel[7]+tmp[6231]*kernel[8];
				ans[6131]<=tmp[6030]*kernel[0]+tmp[6031]*kernel[1]+tmp[6032]*kernel[2]+tmp[6130]*kernel[3]+tmp[6131]*kernel[4]+tmp[6132]*kernel[5]+tmp[6230]*kernel[6]+tmp[6231]*kernel[7]+tmp[6232]*kernel[8];
				ans[6132]<=tmp[6031]*kernel[0]+tmp[6032]*kernel[1]+tmp[6033]*kernel[2]+tmp[6131]*kernel[3]+tmp[6132]*kernel[4]+tmp[6133]*kernel[5]+tmp[6231]*kernel[6]+tmp[6232]*kernel[7]+tmp[6233]*kernel[8];
				ans[6133]<=tmp[6032]*kernel[0]+tmp[6033]*kernel[1]+tmp[6034]*kernel[2]+tmp[6132]*kernel[3]+tmp[6133]*kernel[4]+tmp[6134]*kernel[5]+tmp[6232]*kernel[6]+tmp[6233]*kernel[7]+tmp[6234]*kernel[8];
				ans[6134]<=tmp[6033]*kernel[0]+tmp[6034]*kernel[1]+tmp[6035]*kernel[2]+tmp[6133]*kernel[3]+tmp[6134]*kernel[4]+tmp[6135]*kernel[5]+tmp[6233]*kernel[6]+tmp[6234]*kernel[7]+tmp[6235]*kernel[8];
				ans[6135]<=tmp[6034]*kernel[0]+tmp[6035]*kernel[1]+tmp[6036]*kernel[2]+tmp[6134]*kernel[3]+tmp[6135]*kernel[4]+tmp[6136]*kernel[5]+tmp[6234]*kernel[6]+tmp[6235]*kernel[7]+tmp[6236]*kernel[8];
				ans[6136]<=tmp[6035]*kernel[0]+tmp[6036]*kernel[1]+tmp[6037]*kernel[2]+tmp[6135]*kernel[3]+tmp[6136]*kernel[4]+tmp[6137]*kernel[5]+tmp[6235]*kernel[6]+tmp[6236]*kernel[7]+tmp[6237]*kernel[8];
				ans[6137]<=tmp[6036]*kernel[0]+tmp[6037]*kernel[1]+tmp[6038]*kernel[2]+tmp[6136]*kernel[3]+tmp[6137]*kernel[4]+tmp[6138]*kernel[5]+tmp[6236]*kernel[6]+tmp[6237]*kernel[7]+tmp[6238]*kernel[8];
				ans[6138]<=tmp[6037]*kernel[0]+tmp[6038]*kernel[1]+tmp[6039]*kernel[2]+tmp[6137]*kernel[3]+tmp[6138]*kernel[4]+tmp[6139]*kernel[5]+tmp[6237]*kernel[6]+tmp[6238]*kernel[7]+tmp[6239]*kernel[8];
				ans[6139]<=tmp[6038]*kernel[0]+tmp[6039]*kernel[1]+tmp[6040]*kernel[2]+tmp[6138]*kernel[3]+tmp[6139]*kernel[4]+tmp[6140]*kernel[5]+tmp[6238]*kernel[6]+tmp[6239]*kernel[7]+tmp[6240]*kernel[8];
				ans[6140]<=tmp[6039]*kernel[0]+tmp[6040]*kernel[1]+tmp[6041]*kernel[2]+tmp[6139]*kernel[3]+tmp[6140]*kernel[4]+tmp[6141]*kernel[5]+tmp[6239]*kernel[6]+tmp[6240]*kernel[7]+tmp[6241]*kernel[8];
				ans[6141]<=tmp[6040]*kernel[0]+tmp[6041]*kernel[1]+tmp[6042]*kernel[2]+tmp[6140]*kernel[3]+tmp[6141]*kernel[4]+tmp[6142]*kernel[5]+tmp[6240]*kernel[6]+tmp[6241]*kernel[7]+tmp[6242]*kernel[8];
				ans[6142]<=tmp[6041]*kernel[0]+tmp[6042]*kernel[1]+tmp[6043]*kernel[2]+tmp[6141]*kernel[3]+tmp[6142]*kernel[4]+tmp[6143]*kernel[5]+tmp[6241]*kernel[6]+tmp[6242]*kernel[7]+tmp[6243]*kernel[8];
				ans[6143]<=tmp[6042]*kernel[0]+tmp[6043]*kernel[1]+tmp[6044]*kernel[2]+tmp[6142]*kernel[3]+tmp[6143]*kernel[4]+tmp[6144]*kernel[5]+tmp[6242]*kernel[6]+tmp[6243]*kernel[7]+tmp[6244]*kernel[8];
				ans[6144]<=tmp[6043]*kernel[0]+tmp[6044]*kernel[1]+tmp[6045]*kernel[2]+tmp[6143]*kernel[3]+tmp[6144]*kernel[4]+tmp[6145]*kernel[5]+tmp[6243]*kernel[6]+tmp[6244]*kernel[7]+tmp[6245]*kernel[8];
				ans[6145]<=tmp[6044]*kernel[0]+tmp[6045]*kernel[1]+tmp[6046]*kernel[2]+tmp[6144]*kernel[3]+tmp[6145]*kernel[4]+tmp[6146]*kernel[5]+tmp[6244]*kernel[6]+tmp[6245]*kernel[7]+tmp[6246]*kernel[8];
				ans[6146]<=tmp[6045]*kernel[0]+tmp[6046]*kernel[1]+tmp[6047]*kernel[2]+tmp[6145]*kernel[3]+tmp[6146]*kernel[4]+tmp[6147]*kernel[5]+tmp[6245]*kernel[6]+tmp[6246]*kernel[7]+tmp[6247]*kernel[8];
				ans[6147]<=tmp[6046]*kernel[0]+tmp[6047]*kernel[1]+tmp[6048]*kernel[2]+tmp[6146]*kernel[3]+tmp[6147]*kernel[4]+tmp[6148]*kernel[5]+tmp[6246]*kernel[6]+tmp[6247]*kernel[7]+tmp[6248]*kernel[8];
				ans[6148]<=tmp[6047]*kernel[0]+tmp[6048]*kernel[1]+tmp[6049]*kernel[2]+tmp[6147]*kernel[3]+tmp[6148]*kernel[4]+tmp[6149]*kernel[5]+tmp[6247]*kernel[6]+tmp[6248]*kernel[7]+tmp[6249]*kernel[8];
				ans[6149]<=tmp[6048]*kernel[0]+tmp[6049]*kernel[1]+tmp[6050]*kernel[2]+tmp[6148]*kernel[3]+tmp[6149]*kernel[4]+tmp[6150]*kernel[5]+tmp[6248]*kernel[6]+tmp[6249]*kernel[7]+tmp[6250]*kernel[8];
				ans[6150]<=tmp[6049]*kernel[0]+tmp[6050]*kernel[1]+tmp[6051]*kernel[2]+tmp[6149]*kernel[3]+tmp[6150]*kernel[4]+tmp[6151]*kernel[5]+tmp[6249]*kernel[6]+tmp[6250]*kernel[7]+tmp[6251]*kernel[8];
				ans[6151]<=tmp[6050]*kernel[0]+tmp[6051]*kernel[1]+tmp[6052]*kernel[2]+tmp[6150]*kernel[3]+tmp[6151]*kernel[4]+tmp[6152]*kernel[5]+tmp[6250]*kernel[6]+tmp[6251]*kernel[7]+tmp[6252]*kernel[8];
				ans[6152]<=tmp[6051]*kernel[0]+tmp[6052]*kernel[1]+tmp[6053]*kernel[2]+tmp[6151]*kernel[3]+tmp[6152]*kernel[4]+tmp[6153]*kernel[5]+tmp[6251]*kernel[6]+tmp[6252]*kernel[7]+tmp[6253]*kernel[8];
				ans[6153]<=tmp[6052]*kernel[0]+tmp[6053]*kernel[1]+tmp[6054]*kernel[2]+tmp[6152]*kernel[3]+tmp[6153]*kernel[4]+tmp[6154]*kernel[5]+tmp[6252]*kernel[6]+tmp[6253]*kernel[7]+tmp[6254]*kernel[8];
				ans[6154]<=tmp[6053]*kernel[0]+tmp[6054]*kernel[1]+tmp[6055]*kernel[2]+tmp[6153]*kernel[3]+tmp[6154]*kernel[4]+tmp[6155]*kernel[5]+tmp[6253]*kernel[6]+tmp[6254]*kernel[7]+tmp[6255]*kernel[8];
				ans[6155]<=tmp[6054]*kernel[0]+tmp[6055]*kernel[1]+tmp[6056]*kernel[2]+tmp[6154]*kernel[3]+tmp[6155]*kernel[4]+tmp[6156]*kernel[5]+tmp[6254]*kernel[6]+tmp[6255]*kernel[7]+tmp[6256]*kernel[8];
				ans[6156]<=tmp[6055]*kernel[0]+tmp[6056]*kernel[1]+tmp[6057]*kernel[2]+tmp[6155]*kernel[3]+tmp[6156]*kernel[4]+tmp[6157]*kernel[5]+tmp[6255]*kernel[6]+tmp[6256]*kernel[7]+tmp[6257]*kernel[8];
				ans[6157]<=tmp[6056]*kernel[0]+tmp[6057]*kernel[1]+tmp[6058]*kernel[2]+tmp[6156]*kernel[3]+tmp[6157]*kernel[4]+tmp[6158]*kernel[5]+tmp[6256]*kernel[6]+tmp[6257]*kernel[7]+tmp[6258]*kernel[8];
				ans[6158]<=tmp[6057]*kernel[0]+tmp[6058]*kernel[1]+tmp[6059]*kernel[2]+tmp[6157]*kernel[3]+tmp[6158]*kernel[4]+tmp[6159]*kernel[5]+tmp[6257]*kernel[6]+tmp[6258]*kernel[7]+tmp[6259]*kernel[8];
				ans[6159]<=tmp[6058]*kernel[0]+tmp[6059]*kernel[1]+tmp[6060]*kernel[2]+tmp[6158]*kernel[3]+tmp[6159]*kernel[4]+tmp[6160]*kernel[5]+tmp[6258]*kernel[6]+tmp[6259]*kernel[7]+tmp[6260]*kernel[8];
				ans[6160]<=tmp[6059]*kernel[0]+tmp[6060]*kernel[1]+tmp[6061]*kernel[2]+tmp[6159]*kernel[3]+tmp[6160]*kernel[4]+tmp[6161]*kernel[5]+tmp[6259]*kernel[6]+tmp[6260]*kernel[7]+tmp[6261]*kernel[8];
				ans[6161]<=tmp[6060]*kernel[0]+tmp[6061]*kernel[1]+tmp[6062]*kernel[2]+tmp[6160]*kernel[3]+tmp[6161]*kernel[4]+tmp[6162]*kernel[5]+tmp[6260]*kernel[6]+tmp[6261]*kernel[7]+tmp[6262]*kernel[8];
				ans[6162]<=tmp[6061]*kernel[0]+tmp[6062]*kernel[1]+tmp[6063]*kernel[2]+tmp[6161]*kernel[3]+tmp[6162]*kernel[4]+tmp[6163]*kernel[5]+tmp[6261]*kernel[6]+tmp[6262]*kernel[7]+tmp[6263]*kernel[8];
				ans[6163]<=tmp[6062]*kernel[0]+tmp[6063]*kernel[1]+tmp[6064]*kernel[2]+tmp[6162]*kernel[3]+tmp[6163]*kernel[4]+tmp[6164]*kernel[5]+tmp[6262]*kernel[6]+tmp[6263]*kernel[7]+tmp[6264]*kernel[8];
				ans[6164]<=tmp[6063]*kernel[0]+tmp[6064]*kernel[1]+tmp[6065]*kernel[2]+tmp[6163]*kernel[3]+tmp[6164]*kernel[4]+tmp[6165]*kernel[5]+tmp[6263]*kernel[6]+tmp[6264]*kernel[7]+tmp[6265]*kernel[8];
				ans[6165]<=tmp[6064]*kernel[0]+tmp[6065]*kernel[1]+tmp[6066]*kernel[2]+tmp[6164]*kernel[3]+tmp[6165]*kernel[4]+tmp[6166]*kernel[5]+tmp[6264]*kernel[6]+tmp[6265]*kernel[7]+tmp[6266]*kernel[8];
				ans[6166]<=tmp[6065]*kernel[0]+tmp[6066]*kernel[1]+tmp[6067]*kernel[2]+tmp[6165]*kernel[3]+tmp[6166]*kernel[4]+tmp[6167]*kernel[5]+tmp[6265]*kernel[6]+tmp[6266]*kernel[7]+tmp[6267]*kernel[8];
				ans[6167]<=tmp[6066]*kernel[0]+tmp[6067]*kernel[1]+tmp[6068]*kernel[2]+tmp[6166]*kernel[3]+tmp[6167]*kernel[4]+tmp[6168]*kernel[5]+tmp[6266]*kernel[6]+tmp[6267]*kernel[7]+tmp[6268]*kernel[8];
				ans[6168]<=tmp[6067]*kernel[0]+tmp[6068]*kernel[1]+tmp[6069]*kernel[2]+tmp[6167]*kernel[3]+tmp[6168]*kernel[4]+tmp[6169]*kernel[5]+tmp[6267]*kernel[6]+tmp[6268]*kernel[7]+tmp[6269]*kernel[8];
				ans[6169]<=tmp[6068]*kernel[0]+tmp[6069]*kernel[1]+tmp[6070]*kernel[2]+tmp[6168]*kernel[3]+tmp[6169]*kernel[4]+tmp[6170]*kernel[5]+tmp[6268]*kernel[6]+tmp[6269]*kernel[7]+tmp[6270]*kernel[8];
				ans[6170]<=tmp[6069]*kernel[0]+tmp[6070]*kernel[1]+tmp[6071]*kernel[2]+tmp[6169]*kernel[3]+tmp[6170]*kernel[4]+tmp[6171]*kernel[5]+tmp[6269]*kernel[6]+tmp[6270]*kernel[7]+tmp[6271]*kernel[8];
				ans[6171]<=tmp[6070]*kernel[0]+tmp[6071]*kernel[1]+tmp[6072]*kernel[2]+tmp[6170]*kernel[3]+tmp[6171]*kernel[4]+tmp[6172]*kernel[5]+tmp[6270]*kernel[6]+tmp[6271]*kernel[7]+tmp[6272]*kernel[8];
				ans[6172]<=tmp[6071]*kernel[0]+tmp[6072]*kernel[1]+tmp[6073]*kernel[2]+tmp[6171]*kernel[3]+tmp[6172]*kernel[4]+tmp[6173]*kernel[5]+tmp[6271]*kernel[6]+tmp[6272]*kernel[7]+tmp[6273]*kernel[8];
				ans[6173]<=tmp[6072]*kernel[0]+tmp[6073]*kernel[1]+tmp[6074]*kernel[2]+tmp[6172]*kernel[3]+tmp[6173]*kernel[4]+tmp[6174]*kernel[5]+tmp[6272]*kernel[6]+tmp[6273]*kernel[7]+tmp[6274]*kernel[8];
				ans[6174]<=tmp[6073]*kernel[0]+tmp[6074]*kernel[1]+tmp[6075]*kernel[2]+tmp[6173]*kernel[3]+tmp[6174]*kernel[4]+tmp[6175]*kernel[5]+tmp[6273]*kernel[6]+tmp[6274]*kernel[7]+tmp[6275]*kernel[8];
				ans[6175]<=tmp[6074]*kernel[0]+tmp[6075]*kernel[1]+tmp[6076]*kernel[2]+tmp[6174]*kernel[3]+tmp[6175]*kernel[4]+tmp[6176]*kernel[5]+tmp[6274]*kernel[6]+tmp[6275]*kernel[7]+tmp[6276]*kernel[8];
				ans[6176]<=tmp[6075]*kernel[0]+tmp[6076]*kernel[1]+tmp[6077]*kernel[2]+tmp[6175]*kernel[3]+tmp[6176]*kernel[4]+tmp[6177]*kernel[5]+tmp[6275]*kernel[6]+tmp[6276]*kernel[7]+tmp[6277]*kernel[8];
				ans[6177]<=tmp[6076]*kernel[0]+tmp[6077]*kernel[1]+tmp[6078]*kernel[2]+tmp[6176]*kernel[3]+tmp[6177]*kernel[4]+tmp[6178]*kernel[5]+tmp[6276]*kernel[6]+tmp[6277]*kernel[7]+tmp[6278]*kernel[8];
				ans[6178]<=tmp[6077]*kernel[0]+tmp[6078]*kernel[1]+tmp[6079]*kernel[2]+tmp[6177]*kernel[3]+tmp[6178]*kernel[4]+tmp[6179]*kernel[5]+tmp[6277]*kernel[6]+tmp[6278]*kernel[7]+tmp[6279]*kernel[8];
				ans[6179]<=tmp[6078]*kernel[0]+tmp[6079]*kernel[1]+tmp[6080]*kernel[2]+tmp[6178]*kernel[3]+tmp[6179]*kernel[4]+tmp[6180]*kernel[5]+tmp[6278]*kernel[6]+tmp[6279]*kernel[7]+tmp[6280]*kernel[8];
				ans[6180]<=tmp[6079]*kernel[0]+tmp[6080]*kernel[1]+tmp[6081]*kernel[2]+tmp[6179]*kernel[3]+tmp[6180]*kernel[4]+tmp[6181]*kernel[5]+tmp[6279]*kernel[6]+tmp[6280]*kernel[7]+tmp[6281]*kernel[8];
				ans[6181]<=tmp[6080]*kernel[0]+tmp[6081]*kernel[1]+tmp[6082]*kernel[2]+tmp[6180]*kernel[3]+tmp[6181]*kernel[4]+tmp[6182]*kernel[5]+tmp[6280]*kernel[6]+tmp[6281]*kernel[7]+tmp[6282]*kernel[8];
				ans[6182]<=tmp[6081]*kernel[0]+tmp[6082]*kernel[1]+tmp[6083]*kernel[2]+tmp[6181]*kernel[3]+tmp[6182]*kernel[4]+tmp[6183]*kernel[5]+tmp[6281]*kernel[6]+tmp[6282]*kernel[7]+tmp[6283]*kernel[8];
				ans[6183]<=tmp[6082]*kernel[0]+tmp[6083]*kernel[1]+tmp[6084]*kernel[2]+tmp[6182]*kernel[3]+tmp[6183]*kernel[4]+tmp[6184]*kernel[5]+tmp[6282]*kernel[6]+tmp[6283]*kernel[7]+tmp[6284]*kernel[8];
				ans[6184]<=tmp[6083]*kernel[0]+tmp[6084]*kernel[1]+tmp[6085]*kernel[2]+tmp[6183]*kernel[3]+tmp[6184]*kernel[4]+tmp[6185]*kernel[5]+tmp[6283]*kernel[6]+tmp[6284]*kernel[7]+tmp[6285]*kernel[8];
				ans[6185]<=tmp[6084]*kernel[0]+tmp[6085]*kernel[1]+tmp[6086]*kernel[2]+tmp[6184]*kernel[3]+tmp[6185]*kernel[4]+tmp[6186]*kernel[5]+tmp[6284]*kernel[6]+tmp[6285]*kernel[7]+tmp[6286]*kernel[8];
				ans[6186]<=tmp[6085]*kernel[0]+tmp[6086]*kernel[1]+tmp[6087]*kernel[2]+tmp[6185]*kernel[3]+tmp[6186]*kernel[4]+tmp[6187]*kernel[5]+tmp[6285]*kernel[6]+tmp[6286]*kernel[7]+tmp[6287]*kernel[8];
				ans[6187]<=tmp[6086]*kernel[0]+tmp[6087]*kernel[1]+tmp[6088]*kernel[2]+tmp[6186]*kernel[3]+tmp[6187]*kernel[4]+tmp[6188]*kernel[5]+tmp[6286]*kernel[6]+tmp[6287]*kernel[7]+tmp[6288]*kernel[8];
				ans[6188]<=tmp[6087]*kernel[0]+tmp[6088]*kernel[1]+tmp[6089]*kernel[2]+tmp[6187]*kernel[3]+tmp[6188]*kernel[4]+tmp[6189]*kernel[5]+tmp[6287]*kernel[6]+tmp[6288]*kernel[7]+tmp[6289]*kernel[8];
				ans[6189]<=tmp[6088]*kernel[0]+tmp[6089]*kernel[1]+tmp[6090]*kernel[2]+tmp[6188]*kernel[3]+tmp[6189]*kernel[4]+tmp[6190]*kernel[5]+tmp[6288]*kernel[6]+tmp[6289]*kernel[7]+tmp[6290]*kernel[8];
				ans[6190]<=tmp[6089]*kernel[0]+tmp[6090]*kernel[1]+tmp[6091]*kernel[2]+tmp[6189]*kernel[3]+tmp[6190]*kernel[4]+tmp[6191]*kernel[5]+tmp[6289]*kernel[6]+tmp[6290]*kernel[7]+tmp[6291]*kernel[8];
				ans[6191]<=tmp[6090]*kernel[0]+tmp[6091]*kernel[1]+tmp[6092]*kernel[2]+tmp[6190]*kernel[3]+tmp[6191]*kernel[4]+tmp[6192]*kernel[5]+tmp[6290]*kernel[6]+tmp[6291]*kernel[7]+tmp[6292]*kernel[8];
				ans[6192]<=tmp[6091]*kernel[0]+tmp[6092]*kernel[1]+tmp[6093]*kernel[2]+tmp[6191]*kernel[3]+tmp[6192]*kernel[4]+tmp[6193]*kernel[5]+tmp[6291]*kernel[6]+tmp[6292]*kernel[7]+tmp[6293]*kernel[8];
				ans[6193]<=tmp[6092]*kernel[0]+tmp[6093]*kernel[1]+tmp[6094]*kernel[2]+tmp[6192]*kernel[3]+tmp[6193]*kernel[4]+tmp[6194]*kernel[5]+tmp[6292]*kernel[6]+tmp[6293]*kernel[7]+tmp[6294]*kernel[8];
				ans[6194]<=tmp[6093]*kernel[0]+tmp[6094]*kernel[1]+tmp[6095]*kernel[2]+tmp[6193]*kernel[3]+tmp[6194]*kernel[4]+tmp[6195]*kernel[5]+tmp[6293]*kernel[6]+tmp[6294]*kernel[7]+tmp[6295]*kernel[8];
				ans[6195]<=tmp[6094]*kernel[0]+tmp[6095]*kernel[1]+tmp[6096]*kernel[2]+tmp[6194]*kernel[3]+tmp[6195]*kernel[4]+tmp[6196]*kernel[5]+tmp[6294]*kernel[6]+tmp[6295]*kernel[7]+tmp[6296]*kernel[8];
				ans[6196]<=tmp[6095]*kernel[0]+tmp[6096]*kernel[1]+tmp[6097]*kernel[2]+tmp[6195]*kernel[3]+tmp[6196]*kernel[4]+tmp[6197]*kernel[5]+tmp[6295]*kernel[6]+tmp[6296]*kernel[7]+tmp[6297]*kernel[8];
				ans[6197]<=tmp[6096]*kernel[0]+tmp[6097]*kernel[1]+tmp[6098]*kernel[2]+tmp[6196]*kernel[3]+tmp[6197]*kernel[4]+tmp[6198]*kernel[5]+tmp[6296]*kernel[6]+tmp[6297]*kernel[7]+tmp[6298]*kernel[8];
				ans[6198]<=tmp[6097]*kernel[0]+tmp[6098]*kernel[1]+tmp[6099]*kernel[2]+tmp[6197]*kernel[3]+tmp[6198]*kernel[4]+tmp[6199]*kernel[5]+tmp[6297]*kernel[6]+tmp[6298]*kernel[7]+tmp[6299]*kernel[8];
				ans[6199]<=tmp[6098]*kernel[0]+tmp[6099]*kernel[1]+tmp[6198]*kernel[3]+tmp[6199]*kernel[4]+tmp[6298]*kernel[6]+tmp[6299]*kernel[7];
				ans[6200]<=tmp[6100]*kernel[1]+tmp[6101]*kernel[2]+tmp[6200]*kernel[4]+tmp[6201]*kernel[5]+tmp[6300]*kernel[7]+tmp[6301]*kernel[8];
				ans[6201]<=tmp[6100]*kernel[0]+tmp[6101]*kernel[1]+tmp[6102]*kernel[2]+tmp[6200]*kernel[3]+tmp[6201]*kernel[4]+tmp[6202]*kernel[5]+tmp[6300]*kernel[6]+tmp[6301]*kernel[7]+tmp[6302]*kernel[8];
				ans[6202]<=tmp[6101]*kernel[0]+tmp[6102]*kernel[1]+tmp[6103]*kernel[2]+tmp[6201]*kernel[3]+tmp[6202]*kernel[4]+tmp[6203]*kernel[5]+tmp[6301]*kernel[6]+tmp[6302]*kernel[7]+tmp[6303]*kernel[8];
				ans[6203]<=tmp[6102]*kernel[0]+tmp[6103]*kernel[1]+tmp[6104]*kernel[2]+tmp[6202]*kernel[3]+tmp[6203]*kernel[4]+tmp[6204]*kernel[5]+tmp[6302]*kernel[6]+tmp[6303]*kernel[7]+tmp[6304]*kernel[8];
				ans[6204]<=tmp[6103]*kernel[0]+tmp[6104]*kernel[1]+tmp[6105]*kernel[2]+tmp[6203]*kernel[3]+tmp[6204]*kernel[4]+tmp[6205]*kernel[5]+tmp[6303]*kernel[6]+tmp[6304]*kernel[7]+tmp[6305]*kernel[8];
				ans[6205]<=tmp[6104]*kernel[0]+tmp[6105]*kernel[1]+tmp[6106]*kernel[2]+tmp[6204]*kernel[3]+tmp[6205]*kernel[4]+tmp[6206]*kernel[5]+tmp[6304]*kernel[6]+tmp[6305]*kernel[7]+tmp[6306]*kernel[8];
				ans[6206]<=tmp[6105]*kernel[0]+tmp[6106]*kernel[1]+tmp[6107]*kernel[2]+tmp[6205]*kernel[3]+tmp[6206]*kernel[4]+tmp[6207]*kernel[5]+tmp[6305]*kernel[6]+tmp[6306]*kernel[7]+tmp[6307]*kernel[8];
				ans[6207]<=tmp[6106]*kernel[0]+tmp[6107]*kernel[1]+tmp[6108]*kernel[2]+tmp[6206]*kernel[3]+tmp[6207]*kernel[4]+tmp[6208]*kernel[5]+tmp[6306]*kernel[6]+tmp[6307]*kernel[7]+tmp[6308]*kernel[8];
				ans[6208]<=tmp[6107]*kernel[0]+tmp[6108]*kernel[1]+tmp[6109]*kernel[2]+tmp[6207]*kernel[3]+tmp[6208]*kernel[4]+tmp[6209]*kernel[5]+tmp[6307]*kernel[6]+tmp[6308]*kernel[7]+tmp[6309]*kernel[8];
				ans[6209]<=tmp[6108]*kernel[0]+tmp[6109]*kernel[1]+tmp[6110]*kernel[2]+tmp[6208]*kernel[3]+tmp[6209]*kernel[4]+tmp[6210]*kernel[5]+tmp[6308]*kernel[6]+tmp[6309]*kernel[7]+tmp[6310]*kernel[8];
				ans[6210]<=tmp[6109]*kernel[0]+tmp[6110]*kernel[1]+tmp[6111]*kernel[2]+tmp[6209]*kernel[3]+tmp[6210]*kernel[4]+tmp[6211]*kernel[5]+tmp[6309]*kernel[6]+tmp[6310]*kernel[7]+tmp[6311]*kernel[8];
				ans[6211]<=tmp[6110]*kernel[0]+tmp[6111]*kernel[1]+tmp[6112]*kernel[2]+tmp[6210]*kernel[3]+tmp[6211]*kernel[4]+tmp[6212]*kernel[5]+tmp[6310]*kernel[6]+tmp[6311]*kernel[7]+tmp[6312]*kernel[8];
				ans[6212]<=tmp[6111]*kernel[0]+tmp[6112]*kernel[1]+tmp[6113]*kernel[2]+tmp[6211]*kernel[3]+tmp[6212]*kernel[4]+tmp[6213]*kernel[5]+tmp[6311]*kernel[6]+tmp[6312]*kernel[7]+tmp[6313]*kernel[8];
				ans[6213]<=tmp[6112]*kernel[0]+tmp[6113]*kernel[1]+tmp[6114]*kernel[2]+tmp[6212]*kernel[3]+tmp[6213]*kernel[4]+tmp[6214]*kernel[5]+tmp[6312]*kernel[6]+tmp[6313]*kernel[7]+tmp[6314]*kernel[8];
				ans[6214]<=tmp[6113]*kernel[0]+tmp[6114]*kernel[1]+tmp[6115]*kernel[2]+tmp[6213]*kernel[3]+tmp[6214]*kernel[4]+tmp[6215]*kernel[5]+tmp[6313]*kernel[6]+tmp[6314]*kernel[7]+tmp[6315]*kernel[8];
				ans[6215]<=tmp[6114]*kernel[0]+tmp[6115]*kernel[1]+tmp[6116]*kernel[2]+tmp[6214]*kernel[3]+tmp[6215]*kernel[4]+tmp[6216]*kernel[5]+tmp[6314]*kernel[6]+tmp[6315]*kernel[7]+tmp[6316]*kernel[8];
				ans[6216]<=tmp[6115]*kernel[0]+tmp[6116]*kernel[1]+tmp[6117]*kernel[2]+tmp[6215]*kernel[3]+tmp[6216]*kernel[4]+tmp[6217]*kernel[5]+tmp[6315]*kernel[6]+tmp[6316]*kernel[7]+tmp[6317]*kernel[8];
				ans[6217]<=tmp[6116]*kernel[0]+tmp[6117]*kernel[1]+tmp[6118]*kernel[2]+tmp[6216]*kernel[3]+tmp[6217]*kernel[4]+tmp[6218]*kernel[5]+tmp[6316]*kernel[6]+tmp[6317]*kernel[7]+tmp[6318]*kernel[8];
				ans[6218]<=tmp[6117]*kernel[0]+tmp[6118]*kernel[1]+tmp[6119]*kernel[2]+tmp[6217]*kernel[3]+tmp[6218]*kernel[4]+tmp[6219]*kernel[5]+tmp[6317]*kernel[6]+tmp[6318]*kernel[7]+tmp[6319]*kernel[8];
				ans[6219]<=tmp[6118]*kernel[0]+tmp[6119]*kernel[1]+tmp[6120]*kernel[2]+tmp[6218]*kernel[3]+tmp[6219]*kernel[4]+tmp[6220]*kernel[5]+tmp[6318]*kernel[6]+tmp[6319]*kernel[7]+tmp[6320]*kernel[8];
				ans[6220]<=tmp[6119]*kernel[0]+tmp[6120]*kernel[1]+tmp[6121]*kernel[2]+tmp[6219]*kernel[3]+tmp[6220]*kernel[4]+tmp[6221]*kernel[5]+tmp[6319]*kernel[6]+tmp[6320]*kernel[7]+tmp[6321]*kernel[8];
				ans[6221]<=tmp[6120]*kernel[0]+tmp[6121]*kernel[1]+tmp[6122]*kernel[2]+tmp[6220]*kernel[3]+tmp[6221]*kernel[4]+tmp[6222]*kernel[5]+tmp[6320]*kernel[6]+tmp[6321]*kernel[7]+tmp[6322]*kernel[8];
				ans[6222]<=tmp[6121]*kernel[0]+tmp[6122]*kernel[1]+tmp[6123]*kernel[2]+tmp[6221]*kernel[3]+tmp[6222]*kernel[4]+tmp[6223]*kernel[5]+tmp[6321]*kernel[6]+tmp[6322]*kernel[7]+tmp[6323]*kernel[8];
				ans[6223]<=tmp[6122]*kernel[0]+tmp[6123]*kernel[1]+tmp[6124]*kernel[2]+tmp[6222]*kernel[3]+tmp[6223]*kernel[4]+tmp[6224]*kernel[5]+tmp[6322]*kernel[6]+tmp[6323]*kernel[7]+tmp[6324]*kernel[8];
				ans[6224]<=tmp[6123]*kernel[0]+tmp[6124]*kernel[1]+tmp[6125]*kernel[2]+tmp[6223]*kernel[3]+tmp[6224]*kernel[4]+tmp[6225]*kernel[5]+tmp[6323]*kernel[6]+tmp[6324]*kernel[7]+tmp[6325]*kernel[8];
				ans[6225]<=tmp[6124]*kernel[0]+tmp[6125]*kernel[1]+tmp[6126]*kernel[2]+tmp[6224]*kernel[3]+tmp[6225]*kernel[4]+tmp[6226]*kernel[5]+tmp[6324]*kernel[6]+tmp[6325]*kernel[7]+tmp[6326]*kernel[8];
				ans[6226]<=tmp[6125]*kernel[0]+tmp[6126]*kernel[1]+tmp[6127]*kernel[2]+tmp[6225]*kernel[3]+tmp[6226]*kernel[4]+tmp[6227]*kernel[5]+tmp[6325]*kernel[6]+tmp[6326]*kernel[7]+tmp[6327]*kernel[8];
				ans[6227]<=tmp[6126]*kernel[0]+tmp[6127]*kernel[1]+tmp[6128]*kernel[2]+tmp[6226]*kernel[3]+tmp[6227]*kernel[4]+tmp[6228]*kernel[5]+tmp[6326]*kernel[6]+tmp[6327]*kernel[7]+tmp[6328]*kernel[8];
				ans[6228]<=tmp[6127]*kernel[0]+tmp[6128]*kernel[1]+tmp[6129]*kernel[2]+tmp[6227]*kernel[3]+tmp[6228]*kernel[4]+tmp[6229]*kernel[5]+tmp[6327]*kernel[6]+tmp[6328]*kernel[7]+tmp[6329]*kernel[8];
				ans[6229]<=tmp[6128]*kernel[0]+tmp[6129]*kernel[1]+tmp[6130]*kernel[2]+tmp[6228]*kernel[3]+tmp[6229]*kernel[4]+tmp[6230]*kernel[5]+tmp[6328]*kernel[6]+tmp[6329]*kernel[7]+tmp[6330]*kernel[8];
				ans[6230]<=tmp[6129]*kernel[0]+tmp[6130]*kernel[1]+tmp[6131]*kernel[2]+tmp[6229]*kernel[3]+tmp[6230]*kernel[4]+tmp[6231]*kernel[5]+tmp[6329]*kernel[6]+tmp[6330]*kernel[7]+tmp[6331]*kernel[8];
				ans[6231]<=tmp[6130]*kernel[0]+tmp[6131]*kernel[1]+tmp[6132]*kernel[2]+tmp[6230]*kernel[3]+tmp[6231]*kernel[4]+tmp[6232]*kernel[5]+tmp[6330]*kernel[6]+tmp[6331]*kernel[7]+tmp[6332]*kernel[8];
				ans[6232]<=tmp[6131]*kernel[0]+tmp[6132]*kernel[1]+tmp[6133]*kernel[2]+tmp[6231]*kernel[3]+tmp[6232]*kernel[4]+tmp[6233]*kernel[5]+tmp[6331]*kernel[6]+tmp[6332]*kernel[7]+tmp[6333]*kernel[8];
				ans[6233]<=tmp[6132]*kernel[0]+tmp[6133]*kernel[1]+tmp[6134]*kernel[2]+tmp[6232]*kernel[3]+tmp[6233]*kernel[4]+tmp[6234]*kernel[5]+tmp[6332]*kernel[6]+tmp[6333]*kernel[7]+tmp[6334]*kernel[8];
				ans[6234]<=tmp[6133]*kernel[0]+tmp[6134]*kernel[1]+tmp[6135]*kernel[2]+tmp[6233]*kernel[3]+tmp[6234]*kernel[4]+tmp[6235]*kernel[5]+tmp[6333]*kernel[6]+tmp[6334]*kernel[7]+tmp[6335]*kernel[8];
				ans[6235]<=tmp[6134]*kernel[0]+tmp[6135]*kernel[1]+tmp[6136]*kernel[2]+tmp[6234]*kernel[3]+tmp[6235]*kernel[4]+tmp[6236]*kernel[5]+tmp[6334]*kernel[6]+tmp[6335]*kernel[7]+tmp[6336]*kernel[8];
				ans[6236]<=tmp[6135]*kernel[0]+tmp[6136]*kernel[1]+tmp[6137]*kernel[2]+tmp[6235]*kernel[3]+tmp[6236]*kernel[4]+tmp[6237]*kernel[5]+tmp[6335]*kernel[6]+tmp[6336]*kernel[7]+tmp[6337]*kernel[8];
				ans[6237]<=tmp[6136]*kernel[0]+tmp[6137]*kernel[1]+tmp[6138]*kernel[2]+tmp[6236]*kernel[3]+tmp[6237]*kernel[4]+tmp[6238]*kernel[5]+tmp[6336]*kernel[6]+tmp[6337]*kernel[7]+tmp[6338]*kernel[8];
				ans[6238]<=tmp[6137]*kernel[0]+tmp[6138]*kernel[1]+tmp[6139]*kernel[2]+tmp[6237]*kernel[3]+tmp[6238]*kernel[4]+tmp[6239]*kernel[5]+tmp[6337]*kernel[6]+tmp[6338]*kernel[7]+tmp[6339]*kernel[8];
				ans[6239]<=tmp[6138]*kernel[0]+tmp[6139]*kernel[1]+tmp[6140]*kernel[2]+tmp[6238]*kernel[3]+tmp[6239]*kernel[4]+tmp[6240]*kernel[5]+tmp[6338]*kernel[6]+tmp[6339]*kernel[7]+tmp[6340]*kernel[8];
				ans[6240]<=tmp[6139]*kernel[0]+tmp[6140]*kernel[1]+tmp[6141]*kernel[2]+tmp[6239]*kernel[3]+tmp[6240]*kernel[4]+tmp[6241]*kernel[5]+tmp[6339]*kernel[6]+tmp[6340]*kernel[7]+tmp[6341]*kernel[8];
				ans[6241]<=tmp[6140]*kernel[0]+tmp[6141]*kernel[1]+tmp[6142]*kernel[2]+tmp[6240]*kernel[3]+tmp[6241]*kernel[4]+tmp[6242]*kernel[5]+tmp[6340]*kernel[6]+tmp[6341]*kernel[7]+tmp[6342]*kernel[8];
				ans[6242]<=tmp[6141]*kernel[0]+tmp[6142]*kernel[1]+tmp[6143]*kernel[2]+tmp[6241]*kernel[3]+tmp[6242]*kernel[4]+tmp[6243]*kernel[5]+tmp[6341]*kernel[6]+tmp[6342]*kernel[7]+tmp[6343]*kernel[8];
				ans[6243]<=tmp[6142]*kernel[0]+tmp[6143]*kernel[1]+tmp[6144]*kernel[2]+tmp[6242]*kernel[3]+tmp[6243]*kernel[4]+tmp[6244]*kernel[5]+tmp[6342]*kernel[6]+tmp[6343]*kernel[7]+tmp[6344]*kernel[8];
				ans[6244]<=tmp[6143]*kernel[0]+tmp[6144]*kernel[1]+tmp[6145]*kernel[2]+tmp[6243]*kernel[3]+tmp[6244]*kernel[4]+tmp[6245]*kernel[5]+tmp[6343]*kernel[6]+tmp[6344]*kernel[7]+tmp[6345]*kernel[8];
				ans[6245]<=tmp[6144]*kernel[0]+tmp[6145]*kernel[1]+tmp[6146]*kernel[2]+tmp[6244]*kernel[3]+tmp[6245]*kernel[4]+tmp[6246]*kernel[5]+tmp[6344]*kernel[6]+tmp[6345]*kernel[7]+tmp[6346]*kernel[8];
				ans[6246]<=tmp[6145]*kernel[0]+tmp[6146]*kernel[1]+tmp[6147]*kernel[2]+tmp[6245]*kernel[3]+tmp[6246]*kernel[4]+tmp[6247]*kernel[5]+tmp[6345]*kernel[6]+tmp[6346]*kernel[7]+tmp[6347]*kernel[8];
				ans[6247]<=tmp[6146]*kernel[0]+tmp[6147]*kernel[1]+tmp[6148]*kernel[2]+tmp[6246]*kernel[3]+tmp[6247]*kernel[4]+tmp[6248]*kernel[5]+tmp[6346]*kernel[6]+tmp[6347]*kernel[7]+tmp[6348]*kernel[8];
				ans[6248]<=tmp[6147]*kernel[0]+tmp[6148]*kernel[1]+tmp[6149]*kernel[2]+tmp[6247]*kernel[3]+tmp[6248]*kernel[4]+tmp[6249]*kernel[5]+tmp[6347]*kernel[6]+tmp[6348]*kernel[7]+tmp[6349]*kernel[8];
				ans[6249]<=tmp[6148]*kernel[0]+tmp[6149]*kernel[1]+tmp[6150]*kernel[2]+tmp[6248]*kernel[3]+tmp[6249]*kernel[4]+tmp[6250]*kernel[5]+tmp[6348]*kernel[6]+tmp[6349]*kernel[7]+tmp[6350]*kernel[8];
				ans[6250]<=tmp[6149]*kernel[0]+tmp[6150]*kernel[1]+tmp[6151]*kernel[2]+tmp[6249]*kernel[3]+tmp[6250]*kernel[4]+tmp[6251]*kernel[5]+tmp[6349]*kernel[6]+tmp[6350]*kernel[7]+tmp[6351]*kernel[8];
				ans[6251]<=tmp[6150]*kernel[0]+tmp[6151]*kernel[1]+tmp[6152]*kernel[2]+tmp[6250]*kernel[3]+tmp[6251]*kernel[4]+tmp[6252]*kernel[5]+tmp[6350]*kernel[6]+tmp[6351]*kernel[7]+tmp[6352]*kernel[8];
				ans[6252]<=tmp[6151]*kernel[0]+tmp[6152]*kernel[1]+tmp[6153]*kernel[2]+tmp[6251]*kernel[3]+tmp[6252]*kernel[4]+tmp[6253]*kernel[5]+tmp[6351]*kernel[6]+tmp[6352]*kernel[7]+tmp[6353]*kernel[8];
				ans[6253]<=tmp[6152]*kernel[0]+tmp[6153]*kernel[1]+tmp[6154]*kernel[2]+tmp[6252]*kernel[3]+tmp[6253]*kernel[4]+tmp[6254]*kernel[5]+tmp[6352]*kernel[6]+tmp[6353]*kernel[7]+tmp[6354]*kernel[8];
				ans[6254]<=tmp[6153]*kernel[0]+tmp[6154]*kernel[1]+tmp[6155]*kernel[2]+tmp[6253]*kernel[3]+tmp[6254]*kernel[4]+tmp[6255]*kernel[5]+tmp[6353]*kernel[6]+tmp[6354]*kernel[7]+tmp[6355]*kernel[8];
				ans[6255]<=tmp[6154]*kernel[0]+tmp[6155]*kernel[1]+tmp[6156]*kernel[2]+tmp[6254]*kernel[3]+tmp[6255]*kernel[4]+tmp[6256]*kernel[5]+tmp[6354]*kernel[6]+tmp[6355]*kernel[7]+tmp[6356]*kernel[8];
				ans[6256]<=tmp[6155]*kernel[0]+tmp[6156]*kernel[1]+tmp[6157]*kernel[2]+tmp[6255]*kernel[3]+tmp[6256]*kernel[4]+tmp[6257]*kernel[5]+tmp[6355]*kernel[6]+tmp[6356]*kernel[7]+tmp[6357]*kernel[8];
				ans[6257]<=tmp[6156]*kernel[0]+tmp[6157]*kernel[1]+tmp[6158]*kernel[2]+tmp[6256]*kernel[3]+tmp[6257]*kernel[4]+tmp[6258]*kernel[5]+tmp[6356]*kernel[6]+tmp[6357]*kernel[7]+tmp[6358]*kernel[8];
				ans[6258]<=tmp[6157]*kernel[0]+tmp[6158]*kernel[1]+tmp[6159]*kernel[2]+tmp[6257]*kernel[3]+tmp[6258]*kernel[4]+tmp[6259]*kernel[5]+tmp[6357]*kernel[6]+tmp[6358]*kernel[7]+tmp[6359]*kernel[8];
				ans[6259]<=tmp[6158]*kernel[0]+tmp[6159]*kernel[1]+tmp[6160]*kernel[2]+tmp[6258]*kernel[3]+tmp[6259]*kernel[4]+tmp[6260]*kernel[5]+tmp[6358]*kernel[6]+tmp[6359]*kernel[7]+tmp[6360]*kernel[8];
				ans[6260]<=tmp[6159]*kernel[0]+tmp[6160]*kernel[1]+tmp[6161]*kernel[2]+tmp[6259]*kernel[3]+tmp[6260]*kernel[4]+tmp[6261]*kernel[5]+tmp[6359]*kernel[6]+tmp[6360]*kernel[7]+tmp[6361]*kernel[8];
				ans[6261]<=tmp[6160]*kernel[0]+tmp[6161]*kernel[1]+tmp[6162]*kernel[2]+tmp[6260]*kernel[3]+tmp[6261]*kernel[4]+tmp[6262]*kernel[5]+tmp[6360]*kernel[6]+tmp[6361]*kernel[7]+tmp[6362]*kernel[8];
				ans[6262]<=tmp[6161]*kernel[0]+tmp[6162]*kernel[1]+tmp[6163]*kernel[2]+tmp[6261]*kernel[3]+tmp[6262]*kernel[4]+tmp[6263]*kernel[5]+tmp[6361]*kernel[6]+tmp[6362]*kernel[7]+tmp[6363]*kernel[8];
				ans[6263]<=tmp[6162]*kernel[0]+tmp[6163]*kernel[1]+tmp[6164]*kernel[2]+tmp[6262]*kernel[3]+tmp[6263]*kernel[4]+tmp[6264]*kernel[5]+tmp[6362]*kernel[6]+tmp[6363]*kernel[7]+tmp[6364]*kernel[8];
				ans[6264]<=tmp[6163]*kernel[0]+tmp[6164]*kernel[1]+tmp[6165]*kernel[2]+tmp[6263]*kernel[3]+tmp[6264]*kernel[4]+tmp[6265]*kernel[5]+tmp[6363]*kernel[6]+tmp[6364]*kernel[7]+tmp[6365]*kernel[8];
				ans[6265]<=tmp[6164]*kernel[0]+tmp[6165]*kernel[1]+tmp[6166]*kernel[2]+tmp[6264]*kernel[3]+tmp[6265]*kernel[4]+tmp[6266]*kernel[5]+tmp[6364]*kernel[6]+tmp[6365]*kernel[7]+tmp[6366]*kernel[8];
				ans[6266]<=tmp[6165]*kernel[0]+tmp[6166]*kernel[1]+tmp[6167]*kernel[2]+tmp[6265]*kernel[3]+tmp[6266]*kernel[4]+tmp[6267]*kernel[5]+tmp[6365]*kernel[6]+tmp[6366]*kernel[7]+tmp[6367]*kernel[8];
				ans[6267]<=tmp[6166]*kernel[0]+tmp[6167]*kernel[1]+tmp[6168]*kernel[2]+tmp[6266]*kernel[3]+tmp[6267]*kernel[4]+tmp[6268]*kernel[5]+tmp[6366]*kernel[6]+tmp[6367]*kernel[7]+tmp[6368]*kernel[8];
				ans[6268]<=tmp[6167]*kernel[0]+tmp[6168]*kernel[1]+tmp[6169]*kernel[2]+tmp[6267]*kernel[3]+tmp[6268]*kernel[4]+tmp[6269]*kernel[5]+tmp[6367]*kernel[6]+tmp[6368]*kernel[7]+tmp[6369]*kernel[8];
				ans[6269]<=tmp[6168]*kernel[0]+tmp[6169]*kernel[1]+tmp[6170]*kernel[2]+tmp[6268]*kernel[3]+tmp[6269]*kernel[4]+tmp[6270]*kernel[5]+tmp[6368]*kernel[6]+tmp[6369]*kernel[7]+tmp[6370]*kernel[8];
				ans[6270]<=tmp[6169]*kernel[0]+tmp[6170]*kernel[1]+tmp[6171]*kernel[2]+tmp[6269]*kernel[3]+tmp[6270]*kernel[4]+tmp[6271]*kernel[5]+tmp[6369]*kernel[6]+tmp[6370]*kernel[7]+tmp[6371]*kernel[8];
				ans[6271]<=tmp[6170]*kernel[0]+tmp[6171]*kernel[1]+tmp[6172]*kernel[2]+tmp[6270]*kernel[3]+tmp[6271]*kernel[4]+tmp[6272]*kernel[5]+tmp[6370]*kernel[6]+tmp[6371]*kernel[7]+tmp[6372]*kernel[8];
				ans[6272]<=tmp[6171]*kernel[0]+tmp[6172]*kernel[1]+tmp[6173]*kernel[2]+tmp[6271]*kernel[3]+tmp[6272]*kernel[4]+tmp[6273]*kernel[5]+tmp[6371]*kernel[6]+tmp[6372]*kernel[7]+tmp[6373]*kernel[8];
				ans[6273]<=tmp[6172]*kernel[0]+tmp[6173]*kernel[1]+tmp[6174]*kernel[2]+tmp[6272]*kernel[3]+tmp[6273]*kernel[4]+tmp[6274]*kernel[5]+tmp[6372]*kernel[6]+tmp[6373]*kernel[7]+tmp[6374]*kernel[8];
				ans[6274]<=tmp[6173]*kernel[0]+tmp[6174]*kernel[1]+tmp[6175]*kernel[2]+tmp[6273]*kernel[3]+tmp[6274]*kernel[4]+tmp[6275]*kernel[5]+tmp[6373]*kernel[6]+tmp[6374]*kernel[7]+tmp[6375]*kernel[8];
				ans[6275]<=tmp[6174]*kernel[0]+tmp[6175]*kernel[1]+tmp[6176]*kernel[2]+tmp[6274]*kernel[3]+tmp[6275]*kernel[4]+tmp[6276]*kernel[5]+tmp[6374]*kernel[6]+tmp[6375]*kernel[7]+tmp[6376]*kernel[8];
				ans[6276]<=tmp[6175]*kernel[0]+tmp[6176]*kernel[1]+tmp[6177]*kernel[2]+tmp[6275]*kernel[3]+tmp[6276]*kernel[4]+tmp[6277]*kernel[5]+tmp[6375]*kernel[6]+tmp[6376]*kernel[7]+tmp[6377]*kernel[8];
				ans[6277]<=tmp[6176]*kernel[0]+tmp[6177]*kernel[1]+tmp[6178]*kernel[2]+tmp[6276]*kernel[3]+tmp[6277]*kernel[4]+tmp[6278]*kernel[5]+tmp[6376]*kernel[6]+tmp[6377]*kernel[7]+tmp[6378]*kernel[8];
				ans[6278]<=tmp[6177]*kernel[0]+tmp[6178]*kernel[1]+tmp[6179]*kernel[2]+tmp[6277]*kernel[3]+tmp[6278]*kernel[4]+tmp[6279]*kernel[5]+tmp[6377]*kernel[6]+tmp[6378]*kernel[7]+tmp[6379]*kernel[8];
				ans[6279]<=tmp[6178]*kernel[0]+tmp[6179]*kernel[1]+tmp[6180]*kernel[2]+tmp[6278]*kernel[3]+tmp[6279]*kernel[4]+tmp[6280]*kernel[5]+tmp[6378]*kernel[6]+tmp[6379]*kernel[7]+tmp[6380]*kernel[8];
				ans[6280]<=tmp[6179]*kernel[0]+tmp[6180]*kernel[1]+tmp[6181]*kernel[2]+tmp[6279]*kernel[3]+tmp[6280]*kernel[4]+tmp[6281]*kernel[5]+tmp[6379]*kernel[6]+tmp[6380]*kernel[7]+tmp[6381]*kernel[8];
				ans[6281]<=tmp[6180]*kernel[0]+tmp[6181]*kernel[1]+tmp[6182]*kernel[2]+tmp[6280]*kernel[3]+tmp[6281]*kernel[4]+tmp[6282]*kernel[5]+tmp[6380]*kernel[6]+tmp[6381]*kernel[7]+tmp[6382]*kernel[8];
				ans[6282]<=tmp[6181]*kernel[0]+tmp[6182]*kernel[1]+tmp[6183]*kernel[2]+tmp[6281]*kernel[3]+tmp[6282]*kernel[4]+tmp[6283]*kernel[5]+tmp[6381]*kernel[6]+tmp[6382]*kernel[7]+tmp[6383]*kernel[8];
				ans[6283]<=tmp[6182]*kernel[0]+tmp[6183]*kernel[1]+tmp[6184]*kernel[2]+tmp[6282]*kernel[3]+tmp[6283]*kernel[4]+tmp[6284]*kernel[5]+tmp[6382]*kernel[6]+tmp[6383]*kernel[7]+tmp[6384]*kernel[8];
				ans[6284]<=tmp[6183]*kernel[0]+tmp[6184]*kernel[1]+tmp[6185]*kernel[2]+tmp[6283]*kernel[3]+tmp[6284]*kernel[4]+tmp[6285]*kernel[5]+tmp[6383]*kernel[6]+tmp[6384]*kernel[7]+tmp[6385]*kernel[8];
				ans[6285]<=tmp[6184]*kernel[0]+tmp[6185]*kernel[1]+tmp[6186]*kernel[2]+tmp[6284]*kernel[3]+tmp[6285]*kernel[4]+tmp[6286]*kernel[5]+tmp[6384]*kernel[6]+tmp[6385]*kernel[7]+tmp[6386]*kernel[8];
				ans[6286]<=tmp[6185]*kernel[0]+tmp[6186]*kernel[1]+tmp[6187]*kernel[2]+tmp[6285]*kernel[3]+tmp[6286]*kernel[4]+tmp[6287]*kernel[5]+tmp[6385]*kernel[6]+tmp[6386]*kernel[7]+tmp[6387]*kernel[8];
				ans[6287]<=tmp[6186]*kernel[0]+tmp[6187]*kernel[1]+tmp[6188]*kernel[2]+tmp[6286]*kernel[3]+tmp[6287]*kernel[4]+tmp[6288]*kernel[5]+tmp[6386]*kernel[6]+tmp[6387]*kernel[7]+tmp[6388]*kernel[8];
				ans[6288]<=tmp[6187]*kernel[0]+tmp[6188]*kernel[1]+tmp[6189]*kernel[2]+tmp[6287]*kernel[3]+tmp[6288]*kernel[4]+tmp[6289]*kernel[5]+tmp[6387]*kernel[6]+tmp[6388]*kernel[7]+tmp[6389]*kernel[8];
				ans[6289]<=tmp[6188]*kernel[0]+tmp[6189]*kernel[1]+tmp[6190]*kernel[2]+tmp[6288]*kernel[3]+tmp[6289]*kernel[4]+tmp[6290]*kernel[5]+tmp[6388]*kernel[6]+tmp[6389]*kernel[7]+tmp[6390]*kernel[8];
				ans[6290]<=tmp[6189]*kernel[0]+tmp[6190]*kernel[1]+tmp[6191]*kernel[2]+tmp[6289]*kernel[3]+tmp[6290]*kernel[4]+tmp[6291]*kernel[5]+tmp[6389]*kernel[6]+tmp[6390]*kernel[7]+tmp[6391]*kernel[8];
				ans[6291]<=tmp[6190]*kernel[0]+tmp[6191]*kernel[1]+tmp[6192]*kernel[2]+tmp[6290]*kernel[3]+tmp[6291]*kernel[4]+tmp[6292]*kernel[5]+tmp[6390]*kernel[6]+tmp[6391]*kernel[7]+tmp[6392]*kernel[8];
				ans[6292]<=tmp[6191]*kernel[0]+tmp[6192]*kernel[1]+tmp[6193]*kernel[2]+tmp[6291]*kernel[3]+tmp[6292]*kernel[4]+tmp[6293]*kernel[5]+tmp[6391]*kernel[6]+tmp[6392]*kernel[7]+tmp[6393]*kernel[8];
				ans[6293]<=tmp[6192]*kernel[0]+tmp[6193]*kernel[1]+tmp[6194]*kernel[2]+tmp[6292]*kernel[3]+tmp[6293]*kernel[4]+tmp[6294]*kernel[5]+tmp[6392]*kernel[6]+tmp[6393]*kernel[7]+tmp[6394]*kernel[8];
				ans[6294]<=tmp[6193]*kernel[0]+tmp[6194]*kernel[1]+tmp[6195]*kernel[2]+tmp[6293]*kernel[3]+tmp[6294]*kernel[4]+tmp[6295]*kernel[5]+tmp[6393]*kernel[6]+tmp[6394]*kernel[7]+tmp[6395]*kernel[8];
				ans[6295]<=tmp[6194]*kernel[0]+tmp[6195]*kernel[1]+tmp[6196]*kernel[2]+tmp[6294]*kernel[3]+tmp[6295]*kernel[4]+tmp[6296]*kernel[5]+tmp[6394]*kernel[6]+tmp[6395]*kernel[7]+tmp[6396]*kernel[8];
				ans[6296]<=tmp[6195]*kernel[0]+tmp[6196]*kernel[1]+tmp[6197]*kernel[2]+tmp[6295]*kernel[3]+tmp[6296]*kernel[4]+tmp[6297]*kernel[5]+tmp[6395]*kernel[6]+tmp[6396]*kernel[7]+tmp[6397]*kernel[8];
				ans[6297]<=tmp[6196]*kernel[0]+tmp[6197]*kernel[1]+tmp[6198]*kernel[2]+tmp[6296]*kernel[3]+tmp[6297]*kernel[4]+tmp[6298]*kernel[5]+tmp[6396]*kernel[6]+tmp[6397]*kernel[7]+tmp[6398]*kernel[8];
				ans[6298]<=tmp[6197]*kernel[0]+tmp[6198]*kernel[1]+tmp[6199]*kernel[2]+tmp[6297]*kernel[3]+tmp[6298]*kernel[4]+tmp[6299]*kernel[5]+tmp[6397]*kernel[6]+tmp[6398]*kernel[7]+tmp[6399]*kernel[8];
				ans[6299]<=tmp[6198]*kernel[0]+tmp[6199]*kernel[1]+tmp[6298]*kernel[3]+tmp[6299]*kernel[4]+tmp[6398]*kernel[6]+tmp[6399]*kernel[7];
				ans[6300]<=tmp[6200]*kernel[1]+tmp[6201]*kernel[2]+tmp[6300]*kernel[4]+tmp[6301]*kernel[5]+tmp[6400]*kernel[7]+tmp[6401]*kernel[8];
				ans[6301]<=tmp[6200]*kernel[0]+tmp[6201]*kernel[1]+tmp[6202]*kernel[2]+tmp[6300]*kernel[3]+tmp[6301]*kernel[4]+tmp[6302]*kernel[5]+tmp[6400]*kernel[6]+tmp[6401]*kernel[7]+tmp[6402]*kernel[8];
				ans[6302]<=tmp[6201]*kernel[0]+tmp[6202]*kernel[1]+tmp[6203]*kernel[2]+tmp[6301]*kernel[3]+tmp[6302]*kernel[4]+tmp[6303]*kernel[5]+tmp[6401]*kernel[6]+tmp[6402]*kernel[7]+tmp[6403]*kernel[8];
				ans[6303]<=tmp[6202]*kernel[0]+tmp[6203]*kernel[1]+tmp[6204]*kernel[2]+tmp[6302]*kernel[3]+tmp[6303]*kernel[4]+tmp[6304]*kernel[5]+tmp[6402]*kernel[6]+tmp[6403]*kernel[7]+tmp[6404]*kernel[8];
				ans[6304]<=tmp[6203]*kernel[0]+tmp[6204]*kernel[1]+tmp[6205]*kernel[2]+tmp[6303]*kernel[3]+tmp[6304]*kernel[4]+tmp[6305]*kernel[5]+tmp[6403]*kernel[6]+tmp[6404]*kernel[7]+tmp[6405]*kernel[8];
				ans[6305]<=tmp[6204]*kernel[0]+tmp[6205]*kernel[1]+tmp[6206]*kernel[2]+tmp[6304]*kernel[3]+tmp[6305]*kernel[4]+tmp[6306]*kernel[5]+tmp[6404]*kernel[6]+tmp[6405]*kernel[7]+tmp[6406]*kernel[8];
				ans[6306]<=tmp[6205]*kernel[0]+tmp[6206]*kernel[1]+tmp[6207]*kernel[2]+tmp[6305]*kernel[3]+tmp[6306]*kernel[4]+tmp[6307]*kernel[5]+tmp[6405]*kernel[6]+tmp[6406]*kernel[7]+tmp[6407]*kernel[8];
				ans[6307]<=tmp[6206]*kernel[0]+tmp[6207]*kernel[1]+tmp[6208]*kernel[2]+tmp[6306]*kernel[3]+tmp[6307]*kernel[4]+tmp[6308]*kernel[5]+tmp[6406]*kernel[6]+tmp[6407]*kernel[7]+tmp[6408]*kernel[8];
				ans[6308]<=tmp[6207]*kernel[0]+tmp[6208]*kernel[1]+tmp[6209]*kernel[2]+tmp[6307]*kernel[3]+tmp[6308]*kernel[4]+tmp[6309]*kernel[5]+tmp[6407]*kernel[6]+tmp[6408]*kernel[7]+tmp[6409]*kernel[8];
				ans[6309]<=tmp[6208]*kernel[0]+tmp[6209]*kernel[1]+tmp[6210]*kernel[2]+tmp[6308]*kernel[3]+tmp[6309]*kernel[4]+tmp[6310]*kernel[5]+tmp[6408]*kernel[6]+tmp[6409]*kernel[7]+tmp[6410]*kernel[8];
				ans[6310]<=tmp[6209]*kernel[0]+tmp[6210]*kernel[1]+tmp[6211]*kernel[2]+tmp[6309]*kernel[3]+tmp[6310]*kernel[4]+tmp[6311]*kernel[5]+tmp[6409]*kernel[6]+tmp[6410]*kernel[7]+tmp[6411]*kernel[8];
				ans[6311]<=tmp[6210]*kernel[0]+tmp[6211]*kernel[1]+tmp[6212]*kernel[2]+tmp[6310]*kernel[3]+tmp[6311]*kernel[4]+tmp[6312]*kernel[5]+tmp[6410]*kernel[6]+tmp[6411]*kernel[7]+tmp[6412]*kernel[8];
				ans[6312]<=tmp[6211]*kernel[0]+tmp[6212]*kernel[1]+tmp[6213]*kernel[2]+tmp[6311]*kernel[3]+tmp[6312]*kernel[4]+tmp[6313]*kernel[5]+tmp[6411]*kernel[6]+tmp[6412]*kernel[7]+tmp[6413]*kernel[8];
				ans[6313]<=tmp[6212]*kernel[0]+tmp[6213]*kernel[1]+tmp[6214]*kernel[2]+tmp[6312]*kernel[3]+tmp[6313]*kernel[4]+tmp[6314]*kernel[5]+tmp[6412]*kernel[6]+tmp[6413]*kernel[7]+tmp[6414]*kernel[8];
				ans[6314]<=tmp[6213]*kernel[0]+tmp[6214]*kernel[1]+tmp[6215]*kernel[2]+tmp[6313]*kernel[3]+tmp[6314]*kernel[4]+tmp[6315]*kernel[5]+tmp[6413]*kernel[6]+tmp[6414]*kernel[7]+tmp[6415]*kernel[8];
				ans[6315]<=tmp[6214]*kernel[0]+tmp[6215]*kernel[1]+tmp[6216]*kernel[2]+tmp[6314]*kernel[3]+tmp[6315]*kernel[4]+tmp[6316]*kernel[5]+tmp[6414]*kernel[6]+tmp[6415]*kernel[7]+tmp[6416]*kernel[8];
				ans[6316]<=tmp[6215]*kernel[0]+tmp[6216]*kernel[1]+tmp[6217]*kernel[2]+tmp[6315]*kernel[3]+tmp[6316]*kernel[4]+tmp[6317]*kernel[5]+tmp[6415]*kernel[6]+tmp[6416]*kernel[7]+tmp[6417]*kernel[8];
				ans[6317]<=tmp[6216]*kernel[0]+tmp[6217]*kernel[1]+tmp[6218]*kernel[2]+tmp[6316]*kernel[3]+tmp[6317]*kernel[4]+tmp[6318]*kernel[5]+tmp[6416]*kernel[6]+tmp[6417]*kernel[7]+tmp[6418]*kernel[8];
				ans[6318]<=tmp[6217]*kernel[0]+tmp[6218]*kernel[1]+tmp[6219]*kernel[2]+tmp[6317]*kernel[3]+tmp[6318]*kernel[4]+tmp[6319]*kernel[5]+tmp[6417]*kernel[6]+tmp[6418]*kernel[7]+tmp[6419]*kernel[8];
				ans[6319]<=tmp[6218]*kernel[0]+tmp[6219]*kernel[1]+tmp[6220]*kernel[2]+tmp[6318]*kernel[3]+tmp[6319]*kernel[4]+tmp[6320]*kernel[5]+tmp[6418]*kernel[6]+tmp[6419]*kernel[7]+tmp[6420]*kernel[8];
				ans[6320]<=tmp[6219]*kernel[0]+tmp[6220]*kernel[1]+tmp[6221]*kernel[2]+tmp[6319]*kernel[3]+tmp[6320]*kernel[4]+tmp[6321]*kernel[5]+tmp[6419]*kernel[6]+tmp[6420]*kernel[7]+tmp[6421]*kernel[8];
				ans[6321]<=tmp[6220]*kernel[0]+tmp[6221]*kernel[1]+tmp[6222]*kernel[2]+tmp[6320]*kernel[3]+tmp[6321]*kernel[4]+tmp[6322]*kernel[5]+tmp[6420]*kernel[6]+tmp[6421]*kernel[7]+tmp[6422]*kernel[8];
				ans[6322]<=tmp[6221]*kernel[0]+tmp[6222]*kernel[1]+tmp[6223]*kernel[2]+tmp[6321]*kernel[3]+tmp[6322]*kernel[4]+tmp[6323]*kernel[5]+tmp[6421]*kernel[6]+tmp[6422]*kernel[7]+tmp[6423]*kernel[8];
				ans[6323]<=tmp[6222]*kernel[0]+tmp[6223]*kernel[1]+tmp[6224]*kernel[2]+tmp[6322]*kernel[3]+tmp[6323]*kernel[4]+tmp[6324]*kernel[5]+tmp[6422]*kernel[6]+tmp[6423]*kernel[7]+tmp[6424]*kernel[8];
				ans[6324]<=tmp[6223]*kernel[0]+tmp[6224]*kernel[1]+tmp[6225]*kernel[2]+tmp[6323]*kernel[3]+tmp[6324]*kernel[4]+tmp[6325]*kernel[5]+tmp[6423]*kernel[6]+tmp[6424]*kernel[7]+tmp[6425]*kernel[8];
				ans[6325]<=tmp[6224]*kernel[0]+tmp[6225]*kernel[1]+tmp[6226]*kernel[2]+tmp[6324]*kernel[3]+tmp[6325]*kernel[4]+tmp[6326]*kernel[5]+tmp[6424]*kernel[6]+tmp[6425]*kernel[7]+tmp[6426]*kernel[8];
				ans[6326]<=tmp[6225]*kernel[0]+tmp[6226]*kernel[1]+tmp[6227]*kernel[2]+tmp[6325]*kernel[3]+tmp[6326]*kernel[4]+tmp[6327]*kernel[5]+tmp[6425]*kernel[6]+tmp[6426]*kernel[7]+tmp[6427]*kernel[8];
				ans[6327]<=tmp[6226]*kernel[0]+tmp[6227]*kernel[1]+tmp[6228]*kernel[2]+tmp[6326]*kernel[3]+tmp[6327]*kernel[4]+tmp[6328]*kernel[5]+tmp[6426]*kernel[6]+tmp[6427]*kernel[7]+tmp[6428]*kernel[8];
				ans[6328]<=tmp[6227]*kernel[0]+tmp[6228]*kernel[1]+tmp[6229]*kernel[2]+tmp[6327]*kernel[3]+tmp[6328]*kernel[4]+tmp[6329]*kernel[5]+tmp[6427]*kernel[6]+tmp[6428]*kernel[7]+tmp[6429]*kernel[8];
				ans[6329]<=tmp[6228]*kernel[0]+tmp[6229]*kernel[1]+tmp[6230]*kernel[2]+tmp[6328]*kernel[3]+tmp[6329]*kernel[4]+tmp[6330]*kernel[5]+tmp[6428]*kernel[6]+tmp[6429]*kernel[7]+tmp[6430]*kernel[8];
				ans[6330]<=tmp[6229]*kernel[0]+tmp[6230]*kernel[1]+tmp[6231]*kernel[2]+tmp[6329]*kernel[3]+tmp[6330]*kernel[4]+tmp[6331]*kernel[5]+tmp[6429]*kernel[6]+tmp[6430]*kernel[7]+tmp[6431]*kernel[8];
				ans[6331]<=tmp[6230]*kernel[0]+tmp[6231]*kernel[1]+tmp[6232]*kernel[2]+tmp[6330]*kernel[3]+tmp[6331]*kernel[4]+tmp[6332]*kernel[5]+tmp[6430]*kernel[6]+tmp[6431]*kernel[7]+tmp[6432]*kernel[8];
				ans[6332]<=tmp[6231]*kernel[0]+tmp[6232]*kernel[1]+tmp[6233]*kernel[2]+tmp[6331]*kernel[3]+tmp[6332]*kernel[4]+tmp[6333]*kernel[5]+tmp[6431]*kernel[6]+tmp[6432]*kernel[7]+tmp[6433]*kernel[8];
				ans[6333]<=tmp[6232]*kernel[0]+tmp[6233]*kernel[1]+tmp[6234]*kernel[2]+tmp[6332]*kernel[3]+tmp[6333]*kernel[4]+tmp[6334]*kernel[5]+tmp[6432]*kernel[6]+tmp[6433]*kernel[7]+tmp[6434]*kernel[8];
				ans[6334]<=tmp[6233]*kernel[0]+tmp[6234]*kernel[1]+tmp[6235]*kernel[2]+tmp[6333]*kernel[3]+tmp[6334]*kernel[4]+tmp[6335]*kernel[5]+tmp[6433]*kernel[6]+tmp[6434]*kernel[7]+tmp[6435]*kernel[8];
				ans[6335]<=tmp[6234]*kernel[0]+tmp[6235]*kernel[1]+tmp[6236]*kernel[2]+tmp[6334]*kernel[3]+tmp[6335]*kernel[4]+tmp[6336]*kernel[5]+tmp[6434]*kernel[6]+tmp[6435]*kernel[7]+tmp[6436]*kernel[8];
				ans[6336]<=tmp[6235]*kernel[0]+tmp[6236]*kernel[1]+tmp[6237]*kernel[2]+tmp[6335]*kernel[3]+tmp[6336]*kernel[4]+tmp[6337]*kernel[5]+tmp[6435]*kernel[6]+tmp[6436]*kernel[7]+tmp[6437]*kernel[8];
				ans[6337]<=tmp[6236]*kernel[0]+tmp[6237]*kernel[1]+tmp[6238]*kernel[2]+tmp[6336]*kernel[3]+tmp[6337]*kernel[4]+tmp[6338]*kernel[5]+tmp[6436]*kernel[6]+tmp[6437]*kernel[7]+tmp[6438]*kernel[8];
				ans[6338]<=tmp[6237]*kernel[0]+tmp[6238]*kernel[1]+tmp[6239]*kernel[2]+tmp[6337]*kernel[3]+tmp[6338]*kernel[4]+tmp[6339]*kernel[5]+tmp[6437]*kernel[6]+tmp[6438]*kernel[7]+tmp[6439]*kernel[8];
				ans[6339]<=tmp[6238]*kernel[0]+tmp[6239]*kernel[1]+tmp[6240]*kernel[2]+tmp[6338]*kernel[3]+tmp[6339]*kernel[4]+tmp[6340]*kernel[5]+tmp[6438]*kernel[6]+tmp[6439]*kernel[7]+tmp[6440]*kernel[8];
				ans[6340]<=tmp[6239]*kernel[0]+tmp[6240]*kernel[1]+tmp[6241]*kernel[2]+tmp[6339]*kernel[3]+tmp[6340]*kernel[4]+tmp[6341]*kernel[5]+tmp[6439]*kernel[6]+tmp[6440]*kernel[7]+tmp[6441]*kernel[8];
				ans[6341]<=tmp[6240]*kernel[0]+tmp[6241]*kernel[1]+tmp[6242]*kernel[2]+tmp[6340]*kernel[3]+tmp[6341]*kernel[4]+tmp[6342]*kernel[5]+tmp[6440]*kernel[6]+tmp[6441]*kernel[7]+tmp[6442]*kernel[8];
				ans[6342]<=tmp[6241]*kernel[0]+tmp[6242]*kernel[1]+tmp[6243]*kernel[2]+tmp[6341]*kernel[3]+tmp[6342]*kernel[4]+tmp[6343]*kernel[5]+tmp[6441]*kernel[6]+tmp[6442]*kernel[7]+tmp[6443]*kernel[8];
				ans[6343]<=tmp[6242]*kernel[0]+tmp[6243]*kernel[1]+tmp[6244]*kernel[2]+tmp[6342]*kernel[3]+tmp[6343]*kernel[4]+tmp[6344]*kernel[5]+tmp[6442]*kernel[6]+tmp[6443]*kernel[7]+tmp[6444]*kernel[8];
				ans[6344]<=tmp[6243]*kernel[0]+tmp[6244]*kernel[1]+tmp[6245]*kernel[2]+tmp[6343]*kernel[3]+tmp[6344]*kernel[4]+tmp[6345]*kernel[5]+tmp[6443]*kernel[6]+tmp[6444]*kernel[7]+tmp[6445]*kernel[8];
				ans[6345]<=tmp[6244]*kernel[0]+tmp[6245]*kernel[1]+tmp[6246]*kernel[2]+tmp[6344]*kernel[3]+tmp[6345]*kernel[4]+tmp[6346]*kernel[5]+tmp[6444]*kernel[6]+tmp[6445]*kernel[7]+tmp[6446]*kernel[8];
				ans[6346]<=tmp[6245]*kernel[0]+tmp[6246]*kernel[1]+tmp[6247]*kernel[2]+tmp[6345]*kernel[3]+tmp[6346]*kernel[4]+tmp[6347]*kernel[5]+tmp[6445]*kernel[6]+tmp[6446]*kernel[7]+tmp[6447]*kernel[8];
				ans[6347]<=tmp[6246]*kernel[0]+tmp[6247]*kernel[1]+tmp[6248]*kernel[2]+tmp[6346]*kernel[3]+tmp[6347]*kernel[4]+tmp[6348]*kernel[5]+tmp[6446]*kernel[6]+tmp[6447]*kernel[7]+tmp[6448]*kernel[8];
				ans[6348]<=tmp[6247]*kernel[0]+tmp[6248]*kernel[1]+tmp[6249]*kernel[2]+tmp[6347]*kernel[3]+tmp[6348]*kernel[4]+tmp[6349]*kernel[5]+tmp[6447]*kernel[6]+tmp[6448]*kernel[7]+tmp[6449]*kernel[8];
				ans[6349]<=tmp[6248]*kernel[0]+tmp[6249]*kernel[1]+tmp[6250]*kernel[2]+tmp[6348]*kernel[3]+tmp[6349]*kernel[4]+tmp[6350]*kernel[5]+tmp[6448]*kernel[6]+tmp[6449]*kernel[7]+tmp[6450]*kernel[8];
				ans[6350]<=tmp[6249]*kernel[0]+tmp[6250]*kernel[1]+tmp[6251]*kernel[2]+tmp[6349]*kernel[3]+tmp[6350]*kernel[4]+tmp[6351]*kernel[5]+tmp[6449]*kernel[6]+tmp[6450]*kernel[7]+tmp[6451]*kernel[8];
				ans[6351]<=tmp[6250]*kernel[0]+tmp[6251]*kernel[1]+tmp[6252]*kernel[2]+tmp[6350]*kernel[3]+tmp[6351]*kernel[4]+tmp[6352]*kernel[5]+tmp[6450]*kernel[6]+tmp[6451]*kernel[7]+tmp[6452]*kernel[8];
				ans[6352]<=tmp[6251]*kernel[0]+tmp[6252]*kernel[1]+tmp[6253]*kernel[2]+tmp[6351]*kernel[3]+tmp[6352]*kernel[4]+tmp[6353]*kernel[5]+tmp[6451]*kernel[6]+tmp[6452]*kernel[7]+tmp[6453]*kernel[8];
				ans[6353]<=tmp[6252]*kernel[0]+tmp[6253]*kernel[1]+tmp[6254]*kernel[2]+tmp[6352]*kernel[3]+tmp[6353]*kernel[4]+tmp[6354]*kernel[5]+tmp[6452]*kernel[6]+tmp[6453]*kernel[7]+tmp[6454]*kernel[8];
				ans[6354]<=tmp[6253]*kernel[0]+tmp[6254]*kernel[1]+tmp[6255]*kernel[2]+tmp[6353]*kernel[3]+tmp[6354]*kernel[4]+tmp[6355]*kernel[5]+tmp[6453]*kernel[6]+tmp[6454]*kernel[7]+tmp[6455]*kernel[8];
				ans[6355]<=tmp[6254]*kernel[0]+tmp[6255]*kernel[1]+tmp[6256]*kernel[2]+tmp[6354]*kernel[3]+tmp[6355]*kernel[4]+tmp[6356]*kernel[5]+tmp[6454]*kernel[6]+tmp[6455]*kernel[7]+tmp[6456]*kernel[8];
				ans[6356]<=tmp[6255]*kernel[0]+tmp[6256]*kernel[1]+tmp[6257]*kernel[2]+tmp[6355]*kernel[3]+tmp[6356]*kernel[4]+tmp[6357]*kernel[5]+tmp[6455]*kernel[6]+tmp[6456]*kernel[7]+tmp[6457]*kernel[8];
				ans[6357]<=tmp[6256]*kernel[0]+tmp[6257]*kernel[1]+tmp[6258]*kernel[2]+tmp[6356]*kernel[3]+tmp[6357]*kernel[4]+tmp[6358]*kernel[5]+tmp[6456]*kernel[6]+tmp[6457]*kernel[7]+tmp[6458]*kernel[8];
				ans[6358]<=tmp[6257]*kernel[0]+tmp[6258]*kernel[1]+tmp[6259]*kernel[2]+tmp[6357]*kernel[3]+tmp[6358]*kernel[4]+tmp[6359]*kernel[5]+tmp[6457]*kernel[6]+tmp[6458]*kernel[7]+tmp[6459]*kernel[8];
				ans[6359]<=tmp[6258]*kernel[0]+tmp[6259]*kernel[1]+tmp[6260]*kernel[2]+tmp[6358]*kernel[3]+tmp[6359]*kernel[4]+tmp[6360]*kernel[5]+tmp[6458]*kernel[6]+tmp[6459]*kernel[7]+tmp[6460]*kernel[8];
				ans[6360]<=tmp[6259]*kernel[0]+tmp[6260]*kernel[1]+tmp[6261]*kernel[2]+tmp[6359]*kernel[3]+tmp[6360]*kernel[4]+tmp[6361]*kernel[5]+tmp[6459]*kernel[6]+tmp[6460]*kernel[7]+tmp[6461]*kernel[8];
				ans[6361]<=tmp[6260]*kernel[0]+tmp[6261]*kernel[1]+tmp[6262]*kernel[2]+tmp[6360]*kernel[3]+tmp[6361]*kernel[4]+tmp[6362]*kernel[5]+tmp[6460]*kernel[6]+tmp[6461]*kernel[7]+tmp[6462]*kernel[8];
				ans[6362]<=tmp[6261]*kernel[0]+tmp[6262]*kernel[1]+tmp[6263]*kernel[2]+tmp[6361]*kernel[3]+tmp[6362]*kernel[4]+tmp[6363]*kernel[5]+tmp[6461]*kernel[6]+tmp[6462]*kernel[7]+tmp[6463]*kernel[8];
				ans[6363]<=tmp[6262]*kernel[0]+tmp[6263]*kernel[1]+tmp[6264]*kernel[2]+tmp[6362]*kernel[3]+tmp[6363]*kernel[4]+tmp[6364]*kernel[5]+tmp[6462]*kernel[6]+tmp[6463]*kernel[7]+tmp[6464]*kernel[8];
				ans[6364]<=tmp[6263]*kernel[0]+tmp[6264]*kernel[1]+tmp[6265]*kernel[2]+tmp[6363]*kernel[3]+tmp[6364]*kernel[4]+tmp[6365]*kernel[5]+tmp[6463]*kernel[6]+tmp[6464]*kernel[7]+tmp[6465]*kernel[8];
				ans[6365]<=tmp[6264]*kernel[0]+tmp[6265]*kernel[1]+tmp[6266]*kernel[2]+tmp[6364]*kernel[3]+tmp[6365]*kernel[4]+tmp[6366]*kernel[5]+tmp[6464]*kernel[6]+tmp[6465]*kernel[7]+tmp[6466]*kernel[8];
				ans[6366]<=tmp[6265]*kernel[0]+tmp[6266]*kernel[1]+tmp[6267]*kernel[2]+tmp[6365]*kernel[3]+tmp[6366]*kernel[4]+tmp[6367]*kernel[5]+tmp[6465]*kernel[6]+tmp[6466]*kernel[7]+tmp[6467]*kernel[8];
				ans[6367]<=tmp[6266]*kernel[0]+tmp[6267]*kernel[1]+tmp[6268]*kernel[2]+tmp[6366]*kernel[3]+tmp[6367]*kernel[4]+tmp[6368]*kernel[5]+tmp[6466]*kernel[6]+tmp[6467]*kernel[7]+tmp[6468]*kernel[8];
				ans[6368]<=tmp[6267]*kernel[0]+tmp[6268]*kernel[1]+tmp[6269]*kernel[2]+tmp[6367]*kernel[3]+tmp[6368]*kernel[4]+tmp[6369]*kernel[5]+tmp[6467]*kernel[6]+tmp[6468]*kernel[7]+tmp[6469]*kernel[8];
				ans[6369]<=tmp[6268]*kernel[0]+tmp[6269]*kernel[1]+tmp[6270]*kernel[2]+tmp[6368]*kernel[3]+tmp[6369]*kernel[4]+tmp[6370]*kernel[5]+tmp[6468]*kernel[6]+tmp[6469]*kernel[7]+tmp[6470]*kernel[8];
				ans[6370]<=tmp[6269]*kernel[0]+tmp[6270]*kernel[1]+tmp[6271]*kernel[2]+tmp[6369]*kernel[3]+tmp[6370]*kernel[4]+tmp[6371]*kernel[5]+tmp[6469]*kernel[6]+tmp[6470]*kernel[7]+tmp[6471]*kernel[8];
				ans[6371]<=tmp[6270]*kernel[0]+tmp[6271]*kernel[1]+tmp[6272]*kernel[2]+tmp[6370]*kernel[3]+tmp[6371]*kernel[4]+tmp[6372]*kernel[5]+tmp[6470]*kernel[6]+tmp[6471]*kernel[7]+tmp[6472]*kernel[8];
				ans[6372]<=tmp[6271]*kernel[0]+tmp[6272]*kernel[1]+tmp[6273]*kernel[2]+tmp[6371]*kernel[3]+tmp[6372]*kernel[4]+tmp[6373]*kernel[5]+tmp[6471]*kernel[6]+tmp[6472]*kernel[7]+tmp[6473]*kernel[8];
				ans[6373]<=tmp[6272]*kernel[0]+tmp[6273]*kernel[1]+tmp[6274]*kernel[2]+tmp[6372]*kernel[3]+tmp[6373]*kernel[4]+tmp[6374]*kernel[5]+tmp[6472]*kernel[6]+tmp[6473]*kernel[7]+tmp[6474]*kernel[8];
				ans[6374]<=tmp[6273]*kernel[0]+tmp[6274]*kernel[1]+tmp[6275]*kernel[2]+tmp[6373]*kernel[3]+tmp[6374]*kernel[4]+tmp[6375]*kernel[5]+tmp[6473]*kernel[6]+tmp[6474]*kernel[7]+tmp[6475]*kernel[8];
				ans[6375]<=tmp[6274]*kernel[0]+tmp[6275]*kernel[1]+tmp[6276]*kernel[2]+tmp[6374]*kernel[3]+tmp[6375]*kernel[4]+tmp[6376]*kernel[5]+tmp[6474]*kernel[6]+tmp[6475]*kernel[7]+tmp[6476]*kernel[8];
				ans[6376]<=tmp[6275]*kernel[0]+tmp[6276]*kernel[1]+tmp[6277]*kernel[2]+tmp[6375]*kernel[3]+tmp[6376]*kernel[4]+tmp[6377]*kernel[5]+tmp[6475]*kernel[6]+tmp[6476]*kernel[7]+tmp[6477]*kernel[8];
				ans[6377]<=tmp[6276]*kernel[0]+tmp[6277]*kernel[1]+tmp[6278]*kernel[2]+tmp[6376]*kernel[3]+tmp[6377]*kernel[4]+tmp[6378]*kernel[5]+tmp[6476]*kernel[6]+tmp[6477]*kernel[7]+tmp[6478]*kernel[8];
				ans[6378]<=tmp[6277]*kernel[0]+tmp[6278]*kernel[1]+tmp[6279]*kernel[2]+tmp[6377]*kernel[3]+tmp[6378]*kernel[4]+tmp[6379]*kernel[5]+tmp[6477]*kernel[6]+tmp[6478]*kernel[7]+tmp[6479]*kernel[8];
				ans[6379]<=tmp[6278]*kernel[0]+tmp[6279]*kernel[1]+tmp[6280]*kernel[2]+tmp[6378]*kernel[3]+tmp[6379]*kernel[4]+tmp[6380]*kernel[5]+tmp[6478]*kernel[6]+tmp[6479]*kernel[7]+tmp[6480]*kernel[8];
				ans[6380]<=tmp[6279]*kernel[0]+tmp[6280]*kernel[1]+tmp[6281]*kernel[2]+tmp[6379]*kernel[3]+tmp[6380]*kernel[4]+tmp[6381]*kernel[5]+tmp[6479]*kernel[6]+tmp[6480]*kernel[7]+tmp[6481]*kernel[8];
				ans[6381]<=tmp[6280]*kernel[0]+tmp[6281]*kernel[1]+tmp[6282]*kernel[2]+tmp[6380]*kernel[3]+tmp[6381]*kernel[4]+tmp[6382]*kernel[5]+tmp[6480]*kernel[6]+tmp[6481]*kernel[7]+tmp[6482]*kernel[8];
				ans[6382]<=tmp[6281]*kernel[0]+tmp[6282]*kernel[1]+tmp[6283]*kernel[2]+tmp[6381]*kernel[3]+tmp[6382]*kernel[4]+tmp[6383]*kernel[5]+tmp[6481]*kernel[6]+tmp[6482]*kernel[7]+tmp[6483]*kernel[8];
				ans[6383]<=tmp[6282]*kernel[0]+tmp[6283]*kernel[1]+tmp[6284]*kernel[2]+tmp[6382]*kernel[3]+tmp[6383]*kernel[4]+tmp[6384]*kernel[5]+tmp[6482]*kernel[6]+tmp[6483]*kernel[7]+tmp[6484]*kernel[8];
				ans[6384]<=tmp[6283]*kernel[0]+tmp[6284]*kernel[1]+tmp[6285]*kernel[2]+tmp[6383]*kernel[3]+tmp[6384]*kernel[4]+tmp[6385]*kernel[5]+tmp[6483]*kernel[6]+tmp[6484]*kernel[7]+tmp[6485]*kernel[8];
				ans[6385]<=tmp[6284]*kernel[0]+tmp[6285]*kernel[1]+tmp[6286]*kernel[2]+tmp[6384]*kernel[3]+tmp[6385]*kernel[4]+tmp[6386]*kernel[5]+tmp[6484]*kernel[6]+tmp[6485]*kernel[7]+tmp[6486]*kernel[8];
				ans[6386]<=tmp[6285]*kernel[0]+tmp[6286]*kernel[1]+tmp[6287]*kernel[2]+tmp[6385]*kernel[3]+tmp[6386]*kernel[4]+tmp[6387]*kernel[5]+tmp[6485]*kernel[6]+tmp[6486]*kernel[7]+tmp[6487]*kernel[8];
				ans[6387]<=tmp[6286]*kernel[0]+tmp[6287]*kernel[1]+tmp[6288]*kernel[2]+tmp[6386]*kernel[3]+tmp[6387]*kernel[4]+tmp[6388]*kernel[5]+tmp[6486]*kernel[6]+tmp[6487]*kernel[7]+tmp[6488]*kernel[8];
				ans[6388]<=tmp[6287]*kernel[0]+tmp[6288]*kernel[1]+tmp[6289]*kernel[2]+tmp[6387]*kernel[3]+tmp[6388]*kernel[4]+tmp[6389]*kernel[5]+tmp[6487]*kernel[6]+tmp[6488]*kernel[7]+tmp[6489]*kernel[8];
				ans[6389]<=tmp[6288]*kernel[0]+tmp[6289]*kernel[1]+tmp[6290]*kernel[2]+tmp[6388]*kernel[3]+tmp[6389]*kernel[4]+tmp[6390]*kernel[5]+tmp[6488]*kernel[6]+tmp[6489]*kernel[7]+tmp[6490]*kernel[8];
				ans[6390]<=tmp[6289]*kernel[0]+tmp[6290]*kernel[1]+tmp[6291]*kernel[2]+tmp[6389]*kernel[3]+tmp[6390]*kernel[4]+tmp[6391]*kernel[5]+tmp[6489]*kernel[6]+tmp[6490]*kernel[7]+tmp[6491]*kernel[8];
				ans[6391]<=tmp[6290]*kernel[0]+tmp[6291]*kernel[1]+tmp[6292]*kernel[2]+tmp[6390]*kernel[3]+tmp[6391]*kernel[4]+tmp[6392]*kernel[5]+tmp[6490]*kernel[6]+tmp[6491]*kernel[7]+tmp[6492]*kernel[8];
				ans[6392]<=tmp[6291]*kernel[0]+tmp[6292]*kernel[1]+tmp[6293]*kernel[2]+tmp[6391]*kernel[3]+tmp[6392]*kernel[4]+tmp[6393]*kernel[5]+tmp[6491]*kernel[6]+tmp[6492]*kernel[7]+tmp[6493]*kernel[8];
				ans[6393]<=tmp[6292]*kernel[0]+tmp[6293]*kernel[1]+tmp[6294]*kernel[2]+tmp[6392]*kernel[3]+tmp[6393]*kernel[4]+tmp[6394]*kernel[5]+tmp[6492]*kernel[6]+tmp[6493]*kernel[7]+tmp[6494]*kernel[8];
				ans[6394]<=tmp[6293]*kernel[0]+tmp[6294]*kernel[1]+tmp[6295]*kernel[2]+tmp[6393]*kernel[3]+tmp[6394]*kernel[4]+tmp[6395]*kernel[5]+tmp[6493]*kernel[6]+tmp[6494]*kernel[7]+tmp[6495]*kernel[8];
				ans[6395]<=tmp[6294]*kernel[0]+tmp[6295]*kernel[1]+tmp[6296]*kernel[2]+tmp[6394]*kernel[3]+tmp[6395]*kernel[4]+tmp[6396]*kernel[5]+tmp[6494]*kernel[6]+tmp[6495]*kernel[7]+tmp[6496]*kernel[8];
				ans[6396]<=tmp[6295]*kernel[0]+tmp[6296]*kernel[1]+tmp[6297]*kernel[2]+tmp[6395]*kernel[3]+tmp[6396]*kernel[4]+tmp[6397]*kernel[5]+tmp[6495]*kernel[6]+tmp[6496]*kernel[7]+tmp[6497]*kernel[8];
				ans[6397]<=tmp[6296]*kernel[0]+tmp[6297]*kernel[1]+tmp[6298]*kernel[2]+tmp[6396]*kernel[3]+tmp[6397]*kernel[4]+tmp[6398]*kernel[5]+tmp[6496]*kernel[6]+tmp[6497]*kernel[7]+tmp[6498]*kernel[8];
				ans[6398]<=tmp[6297]*kernel[0]+tmp[6298]*kernel[1]+tmp[6299]*kernel[2]+tmp[6397]*kernel[3]+tmp[6398]*kernel[4]+tmp[6399]*kernel[5]+tmp[6497]*kernel[6]+tmp[6498]*kernel[7]+tmp[6499]*kernel[8];
				ans[6399]<=tmp[6298]*kernel[0]+tmp[6299]*kernel[1]+tmp[6398]*kernel[3]+tmp[6399]*kernel[4]+tmp[6498]*kernel[6]+tmp[6499]*kernel[7];
				ans[6400]<=tmp[6300]*kernel[1]+tmp[6301]*kernel[2]+tmp[6400]*kernel[4]+tmp[6401]*kernel[5]+tmp[6500]*kernel[7]+tmp[6501]*kernel[8];
				ans[6401]<=tmp[6300]*kernel[0]+tmp[6301]*kernel[1]+tmp[6302]*kernel[2]+tmp[6400]*kernel[3]+tmp[6401]*kernel[4]+tmp[6402]*kernel[5]+tmp[6500]*kernel[6]+tmp[6501]*kernel[7]+tmp[6502]*kernel[8];
				ans[6402]<=tmp[6301]*kernel[0]+tmp[6302]*kernel[1]+tmp[6303]*kernel[2]+tmp[6401]*kernel[3]+tmp[6402]*kernel[4]+tmp[6403]*kernel[5]+tmp[6501]*kernel[6]+tmp[6502]*kernel[7]+tmp[6503]*kernel[8];
				ans[6403]<=tmp[6302]*kernel[0]+tmp[6303]*kernel[1]+tmp[6304]*kernel[2]+tmp[6402]*kernel[3]+tmp[6403]*kernel[4]+tmp[6404]*kernel[5]+tmp[6502]*kernel[6]+tmp[6503]*kernel[7]+tmp[6504]*kernel[8];
				ans[6404]<=tmp[6303]*kernel[0]+tmp[6304]*kernel[1]+tmp[6305]*kernel[2]+tmp[6403]*kernel[3]+tmp[6404]*kernel[4]+tmp[6405]*kernel[5]+tmp[6503]*kernel[6]+tmp[6504]*kernel[7]+tmp[6505]*kernel[8];
				ans[6405]<=tmp[6304]*kernel[0]+tmp[6305]*kernel[1]+tmp[6306]*kernel[2]+tmp[6404]*kernel[3]+tmp[6405]*kernel[4]+tmp[6406]*kernel[5]+tmp[6504]*kernel[6]+tmp[6505]*kernel[7]+tmp[6506]*kernel[8];
				ans[6406]<=tmp[6305]*kernel[0]+tmp[6306]*kernel[1]+tmp[6307]*kernel[2]+tmp[6405]*kernel[3]+tmp[6406]*kernel[4]+tmp[6407]*kernel[5]+tmp[6505]*kernel[6]+tmp[6506]*kernel[7]+tmp[6507]*kernel[8];
				ans[6407]<=tmp[6306]*kernel[0]+tmp[6307]*kernel[1]+tmp[6308]*kernel[2]+tmp[6406]*kernel[3]+tmp[6407]*kernel[4]+tmp[6408]*kernel[5]+tmp[6506]*kernel[6]+tmp[6507]*kernel[7]+tmp[6508]*kernel[8];
				ans[6408]<=tmp[6307]*kernel[0]+tmp[6308]*kernel[1]+tmp[6309]*kernel[2]+tmp[6407]*kernel[3]+tmp[6408]*kernel[4]+tmp[6409]*kernel[5]+tmp[6507]*kernel[6]+tmp[6508]*kernel[7]+tmp[6509]*kernel[8];
				ans[6409]<=tmp[6308]*kernel[0]+tmp[6309]*kernel[1]+tmp[6310]*kernel[2]+tmp[6408]*kernel[3]+tmp[6409]*kernel[4]+tmp[6410]*kernel[5]+tmp[6508]*kernel[6]+tmp[6509]*kernel[7]+tmp[6510]*kernel[8];
				ans[6410]<=tmp[6309]*kernel[0]+tmp[6310]*kernel[1]+tmp[6311]*kernel[2]+tmp[6409]*kernel[3]+tmp[6410]*kernel[4]+tmp[6411]*kernel[5]+tmp[6509]*kernel[6]+tmp[6510]*kernel[7]+tmp[6511]*kernel[8];
				ans[6411]<=tmp[6310]*kernel[0]+tmp[6311]*kernel[1]+tmp[6312]*kernel[2]+tmp[6410]*kernel[3]+tmp[6411]*kernel[4]+tmp[6412]*kernel[5]+tmp[6510]*kernel[6]+tmp[6511]*kernel[7]+tmp[6512]*kernel[8];
				ans[6412]<=tmp[6311]*kernel[0]+tmp[6312]*kernel[1]+tmp[6313]*kernel[2]+tmp[6411]*kernel[3]+tmp[6412]*kernel[4]+tmp[6413]*kernel[5]+tmp[6511]*kernel[6]+tmp[6512]*kernel[7]+tmp[6513]*kernel[8];
				ans[6413]<=tmp[6312]*kernel[0]+tmp[6313]*kernel[1]+tmp[6314]*kernel[2]+tmp[6412]*kernel[3]+tmp[6413]*kernel[4]+tmp[6414]*kernel[5]+tmp[6512]*kernel[6]+tmp[6513]*kernel[7]+tmp[6514]*kernel[8];
				ans[6414]<=tmp[6313]*kernel[0]+tmp[6314]*kernel[1]+tmp[6315]*kernel[2]+tmp[6413]*kernel[3]+tmp[6414]*kernel[4]+tmp[6415]*kernel[5]+tmp[6513]*kernel[6]+tmp[6514]*kernel[7]+tmp[6515]*kernel[8];
				ans[6415]<=tmp[6314]*kernel[0]+tmp[6315]*kernel[1]+tmp[6316]*kernel[2]+tmp[6414]*kernel[3]+tmp[6415]*kernel[4]+tmp[6416]*kernel[5]+tmp[6514]*kernel[6]+tmp[6515]*kernel[7]+tmp[6516]*kernel[8];
				ans[6416]<=tmp[6315]*kernel[0]+tmp[6316]*kernel[1]+tmp[6317]*kernel[2]+tmp[6415]*kernel[3]+tmp[6416]*kernel[4]+tmp[6417]*kernel[5]+tmp[6515]*kernel[6]+tmp[6516]*kernel[7]+tmp[6517]*kernel[8];
				ans[6417]<=tmp[6316]*kernel[0]+tmp[6317]*kernel[1]+tmp[6318]*kernel[2]+tmp[6416]*kernel[3]+tmp[6417]*kernel[4]+tmp[6418]*kernel[5]+tmp[6516]*kernel[6]+tmp[6517]*kernel[7]+tmp[6518]*kernel[8];
				ans[6418]<=tmp[6317]*kernel[0]+tmp[6318]*kernel[1]+tmp[6319]*kernel[2]+tmp[6417]*kernel[3]+tmp[6418]*kernel[4]+tmp[6419]*kernel[5]+tmp[6517]*kernel[6]+tmp[6518]*kernel[7]+tmp[6519]*kernel[8];
				ans[6419]<=tmp[6318]*kernel[0]+tmp[6319]*kernel[1]+tmp[6320]*kernel[2]+tmp[6418]*kernel[3]+tmp[6419]*kernel[4]+tmp[6420]*kernel[5]+tmp[6518]*kernel[6]+tmp[6519]*kernel[7]+tmp[6520]*kernel[8];
				ans[6420]<=tmp[6319]*kernel[0]+tmp[6320]*kernel[1]+tmp[6321]*kernel[2]+tmp[6419]*kernel[3]+tmp[6420]*kernel[4]+tmp[6421]*kernel[5]+tmp[6519]*kernel[6]+tmp[6520]*kernel[7]+tmp[6521]*kernel[8];
				ans[6421]<=tmp[6320]*kernel[0]+tmp[6321]*kernel[1]+tmp[6322]*kernel[2]+tmp[6420]*kernel[3]+tmp[6421]*kernel[4]+tmp[6422]*kernel[5]+tmp[6520]*kernel[6]+tmp[6521]*kernel[7]+tmp[6522]*kernel[8];
				ans[6422]<=tmp[6321]*kernel[0]+tmp[6322]*kernel[1]+tmp[6323]*kernel[2]+tmp[6421]*kernel[3]+tmp[6422]*kernel[4]+tmp[6423]*kernel[5]+tmp[6521]*kernel[6]+tmp[6522]*kernel[7]+tmp[6523]*kernel[8];
				ans[6423]<=tmp[6322]*kernel[0]+tmp[6323]*kernel[1]+tmp[6324]*kernel[2]+tmp[6422]*kernel[3]+tmp[6423]*kernel[4]+tmp[6424]*kernel[5]+tmp[6522]*kernel[6]+tmp[6523]*kernel[7]+tmp[6524]*kernel[8];
				ans[6424]<=tmp[6323]*kernel[0]+tmp[6324]*kernel[1]+tmp[6325]*kernel[2]+tmp[6423]*kernel[3]+tmp[6424]*kernel[4]+tmp[6425]*kernel[5]+tmp[6523]*kernel[6]+tmp[6524]*kernel[7]+tmp[6525]*kernel[8];
				ans[6425]<=tmp[6324]*kernel[0]+tmp[6325]*kernel[1]+tmp[6326]*kernel[2]+tmp[6424]*kernel[3]+tmp[6425]*kernel[4]+tmp[6426]*kernel[5]+tmp[6524]*kernel[6]+tmp[6525]*kernel[7]+tmp[6526]*kernel[8];
				ans[6426]<=tmp[6325]*kernel[0]+tmp[6326]*kernel[1]+tmp[6327]*kernel[2]+tmp[6425]*kernel[3]+tmp[6426]*kernel[4]+tmp[6427]*kernel[5]+tmp[6525]*kernel[6]+tmp[6526]*kernel[7]+tmp[6527]*kernel[8];
				ans[6427]<=tmp[6326]*kernel[0]+tmp[6327]*kernel[1]+tmp[6328]*kernel[2]+tmp[6426]*kernel[3]+tmp[6427]*kernel[4]+tmp[6428]*kernel[5]+tmp[6526]*kernel[6]+tmp[6527]*kernel[7]+tmp[6528]*kernel[8];
				ans[6428]<=tmp[6327]*kernel[0]+tmp[6328]*kernel[1]+tmp[6329]*kernel[2]+tmp[6427]*kernel[3]+tmp[6428]*kernel[4]+tmp[6429]*kernel[5]+tmp[6527]*kernel[6]+tmp[6528]*kernel[7]+tmp[6529]*kernel[8];
				ans[6429]<=tmp[6328]*kernel[0]+tmp[6329]*kernel[1]+tmp[6330]*kernel[2]+tmp[6428]*kernel[3]+tmp[6429]*kernel[4]+tmp[6430]*kernel[5]+tmp[6528]*kernel[6]+tmp[6529]*kernel[7]+tmp[6530]*kernel[8];
				ans[6430]<=tmp[6329]*kernel[0]+tmp[6330]*kernel[1]+tmp[6331]*kernel[2]+tmp[6429]*kernel[3]+tmp[6430]*kernel[4]+tmp[6431]*kernel[5]+tmp[6529]*kernel[6]+tmp[6530]*kernel[7]+tmp[6531]*kernel[8];
				ans[6431]<=tmp[6330]*kernel[0]+tmp[6331]*kernel[1]+tmp[6332]*kernel[2]+tmp[6430]*kernel[3]+tmp[6431]*kernel[4]+tmp[6432]*kernel[5]+tmp[6530]*kernel[6]+tmp[6531]*kernel[7]+tmp[6532]*kernel[8];
				ans[6432]<=tmp[6331]*kernel[0]+tmp[6332]*kernel[1]+tmp[6333]*kernel[2]+tmp[6431]*kernel[3]+tmp[6432]*kernel[4]+tmp[6433]*kernel[5]+tmp[6531]*kernel[6]+tmp[6532]*kernel[7]+tmp[6533]*kernel[8];
				ans[6433]<=tmp[6332]*kernel[0]+tmp[6333]*kernel[1]+tmp[6334]*kernel[2]+tmp[6432]*kernel[3]+tmp[6433]*kernel[4]+tmp[6434]*kernel[5]+tmp[6532]*kernel[6]+tmp[6533]*kernel[7]+tmp[6534]*kernel[8];
				ans[6434]<=tmp[6333]*kernel[0]+tmp[6334]*kernel[1]+tmp[6335]*kernel[2]+tmp[6433]*kernel[3]+tmp[6434]*kernel[4]+tmp[6435]*kernel[5]+tmp[6533]*kernel[6]+tmp[6534]*kernel[7]+tmp[6535]*kernel[8];
				ans[6435]<=tmp[6334]*kernel[0]+tmp[6335]*kernel[1]+tmp[6336]*kernel[2]+tmp[6434]*kernel[3]+tmp[6435]*kernel[4]+tmp[6436]*kernel[5]+tmp[6534]*kernel[6]+tmp[6535]*kernel[7]+tmp[6536]*kernel[8];
				ans[6436]<=tmp[6335]*kernel[0]+tmp[6336]*kernel[1]+tmp[6337]*kernel[2]+tmp[6435]*kernel[3]+tmp[6436]*kernel[4]+tmp[6437]*kernel[5]+tmp[6535]*kernel[6]+tmp[6536]*kernel[7]+tmp[6537]*kernel[8];
				ans[6437]<=tmp[6336]*kernel[0]+tmp[6337]*kernel[1]+tmp[6338]*kernel[2]+tmp[6436]*kernel[3]+tmp[6437]*kernel[4]+tmp[6438]*kernel[5]+tmp[6536]*kernel[6]+tmp[6537]*kernel[7]+tmp[6538]*kernel[8];
				ans[6438]<=tmp[6337]*kernel[0]+tmp[6338]*kernel[1]+tmp[6339]*kernel[2]+tmp[6437]*kernel[3]+tmp[6438]*kernel[4]+tmp[6439]*kernel[5]+tmp[6537]*kernel[6]+tmp[6538]*kernel[7]+tmp[6539]*kernel[8];
				ans[6439]<=tmp[6338]*kernel[0]+tmp[6339]*kernel[1]+tmp[6340]*kernel[2]+tmp[6438]*kernel[3]+tmp[6439]*kernel[4]+tmp[6440]*kernel[5]+tmp[6538]*kernel[6]+tmp[6539]*kernel[7]+tmp[6540]*kernel[8];
				ans[6440]<=tmp[6339]*kernel[0]+tmp[6340]*kernel[1]+tmp[6341]*kernel[2]+tmp[6439]*kernel[3]+tmp[6440]*kernel[4]+tmp[6441]*kernel[5]+tmp[6539]*kernel[6]+tmp[6540]*kernel[7]+tmp[6541]*kernel[8];
				ans[6441]<=tmp[6340]*kernel[0]+tmp[6341]*kernel[1]+tmp[6342]*kernel[2]+tmp[6440]*kernel[3]+tmp[6441]*kernel[4]+tmp[6442]*kernel[5]+tmp[6540]*kernel[6]+tmp[6541]*kernel[7]+tmp[6542]*kernel[8];
				ans[6442]<=tmp[6341]*kernel[0]+tmp[6342]*kernel[1]+tmp[6343]*kernel[2]+tmp[6441]*kernel[3]+tmp[6442]*kernel[4]+tmp[6443]*kernel[5]+tmp[6541]*kernel[6]+tmp[6542]*kernel[7]+tmp[6543]*kernel[8];
				ans[6443]<=tmp[6342]*kernel[0]+tmp[6343]*kernel[1]+tmp[6344]*kernel[2]+tmp[6442]*kernel[3]+tmp[6443]*kernel[4]+tmp[6444]*kernel[5]+tmp[6542]*kernel[6]+tmp[6543]*kernel[7]+tmp[6544]*kernel[8];
				ans[6444]<=tmp[6343]*kernel[0]+tmp[6344]*kernel[1]+tmp[6345]*kernel[2]+tmp[6443]*kernel[3]+tmp[6444]*kernel[4]+tmp[6445]*kernel[5]+tmp[6543]*kernel[6]+tmp[6544]*kernel[7]+tmp[6545]*kernel[8];
				ans[6445]<=tmp[6344]*kernel[0]+tmp[6345]*kernel[1]+tmp[6346]*kernel[2]+tmp[6444]*kernel[3]+tmp[6445]*kernel[4]+tmp[6446]*kernel[5]+tmp[6544]*kernel[6]+tmp[6545]*kernel[7]+tmp[6546]*kernel[8];
				ans[6446]<=tmp[6345]*kernel[0]+tmp[6346]*kernel[1]+tmp[6347]*kernel[2]+tmp[6445]*kernel[3]+tmp[6446]*kernel[4]+tmp[6447]*kernel[5]+tmp[6545]*kernel[6]+tmp[6546]*kernel[7]+tmp[6547]*kernel[8];
				ans[6447]<=tmp[6346]*kernel[0]+tmp[6347]*kernel[1]+tmp[6348]*kernel[2]+tmp[6446]*kernel[3]+tmp[6447]*kernel[4]+tmp[6448]*kernel[5]+tmp[6546]*kernel[6]+tmp[6547]*kernel[7]+tmp[6548]*kernel[8];
				ans[6448]<=tmp[6347]*kernel[0]+tmp[6348]*kernel[1]+tmp[6349]*kernel[2]+tmp[6447]*kernel[3]+tmp[6448]*kernel[4]+tmp[6449]*kernel[5]+tmp[6547]*kernel[6]+tmp[6548]*kernel[7]+tmp[6549]*kernel[8];
				ans[6449]<=tmp[6348]*kernel[0]+tmp[6349]*kernel[1]+tmp[6350]*kernel[2]+tmp[6448]*kernel[3]+tmp[6449]*kernel[4]+tmp[6450]*kernel[5]+tmp[6548]*kernel[6]+tmp[6549]*kernel[7]+tmp[6550]*kernel[8];
				ans[6450]<=tmp[6349]*kernel[0]+tmp[6350]*kernel[1]+tmp[6351]*kernel[2]+tmp[6449]*kernel[3]+tmp[6450]*kernel[4]+tmp[6451]*kernel[5]+tmp[6549]*kernel[6]+tmp[6550]*kernel[7]+tmp[6551]*kernel[8];
				ans[6451]<=tmp[6350]*kernel[0]+tmp[6351]*kernel[1]+tmp[6352]*kernel[2]+tmp[6450]*kernel[3]+tmp[6451]*kernel[4]+tmp[6452]*kernel[5]+tmp[6550]*kernel[6]+tmp[6551]*kernel[7]+tmp[6552]*kernel[8];
				ans[6452]<=tmp[6351]*kernel[0]+tmp[6352]*kernel[1]+tmp[6353]*kernel[2]+tmp[6451]*kernel[3]+tmp[6452]*kernel[4]+tmp[6453]*kernel[5]+tmp[6551]*kernel[6]+tmp[6552]*kernel[7]+tmp[6553]*kernel[8];
				ans[6453]<=tmp[6352]*kernel[0]+tmp[6353]*kernel[1]+tmp[6354]*kernel[2]+tmp[6452]*kernel[3]+tmp[6453]*kernel[4]+tmp[6454]*kernel[5]+tmp[6552]*kernel[6]+tmp[6553]*kernel[7]+tmp[6554]*kernel[8];
				ans[6454]<=tmp[6353]*kernel[0]+tmp[6354]*kernel[1]+tmp[6355]*kernel[2]+tmp[6453]*kernel[3]+tmp[6454]*kernel[4]+tmp[6455]*kernel[5]+tmp[6553]*kernel[6]+tmp[6554]*kernel[7]+tmp[6555]*kernel[8];
				ans[6455]<=tmp[6354]*kernel[0]+tmp[6355]*kernel[1]+tmp[6356]*kernel[2]+tmp[6454]*kernel[3]+tmp[6455]*kernel[4]+tmp[6456]*kernel[5]+tmp[6554]*kernel[6]+tmp[6555]*kernel[7]+tmp[6556]*kernel[8];
				ans[6456]<=tmp[6355]*kernel[0]+tmp[6356]*kernel[1]+tmp[6357]*kernel[2]+tmp[6455]*kernel[3]+tmp[6456]*kernel[4]+tmp[6457]*kernel[5]+tmp[6555]*kernel[6]+tmp[6556]*kernel[7]+tmp[6557]*kernel[8];
				ans[6457]<=tmp[6356]*kernel[0]+tmp[6357]*kernel[1]+tmp[6358]*kernel[2]+tmp[6456]*kernel[3]+tmp[6457]*kernel[4]+tmp[6458]*kernel[5]+tmp[6556]*kernel[6]+tmp[6557]*kernel[7]+tmp[6558]*kernel[8];
				ans[6458]<=tmp[6357]*kernel[0]+tmp[6358]*kernel[1]+tmp[6359]*kernel[2]+tmp[6457]*kernel[3]+tmp[6458]*kernel[4]+tmp[6459]*kernel[5]+tmp[6557]*kernel[6]+tmp[6558]*kernel[7]+tmp[6559]*kernel[8];
				ans[6459]<=tmp[6358]*kernel[0]+tmp[6359]*kernel[1]+tmp[6360]*kernel[2]+tmp[6458]*kernel[3]+tmp[6459]*kernel[4]+tmp[6460]*kernel[5]+tmp[6558]*kernel[6]+tmp[6559]*kernel[7]+tmp[6560]*kernel[8];
				ans[6460]<=tmp[6359]*kernel[0]+tmp[6360]*kernel[1]+tmp[6361]*kernel[2]+tmp[6459]*kernel[3]+tmp[6460]*kernel[4]+tmp[6461]*kernel[5]+tmp[6559]*kernel[6]+tmp[6560]*kernel[7]+tmp[6561]*kernel[8];
				ans[6461]<=tmp[6360]*kernel[0]+tmp[6361]*kernel[1]+tmp[6362]*kernel[2]+tmp[6460]*kernel[3]+tmp[6461]*kernel[4]+tmp[6462]*kernel[5]+tmp[6560]*kernel[6]+tmp[6561]*kernel[7]+tmp[6562]*kernel[8];
				ans[6462]<=tmp[6361]*kernel[0]+tmp[6362]*kernel[1]+tmp[6363]*kernel[2]+tmp[6461]*kernel[3]+tmp[6462]*kernel[4]+tmp[6463]*kernel[5]+tmp[6561]*kernel[6]+tmp[6562]*kernel[7]+tmp[6563]*kernel[8];
				ans[6463]<=tmp[6362]*kernel[0]+tmp[6363]*kernel[1]+tmp[6364]*kernel[2]+tmp[6462]*kernel[3]+tmp[6463]*kernel[4]+tmp[6464]*kernel[5]+tmp[6562]*kernel[6]+tmp[6563]*kernel[7]+tmp[6564]*kernel[8];
				ans[6464]<=tmp[6363]*kernel[0]+tmp[6364]*kernel[1]+tmp[6365]*kernel[2]+tmp[6463]*kernel[3]+tmp[6464]*kernel[4]+tmp[6465]*kernel[5]+tmp[6563]*kernel[6]+tmp[6564]*kernel[7]+tmp[6565]*kernel[8];
				ans[6465]<=tmp[6364]*kernel[0]+tmp[6365]*kernel[1]+tmp[6366]*kernel[2]+tmp[6464]*kernel[3]+tmp[6465]*kernel[4]+tmp[6466]*kernel[5]+tmp[6564]*kernel[6]+tmp[6565]*kernel[7]+tmp[6566]*kernel[8];
				ans[6466]<=tmp[6365]*kernel[0]+tmp[6366]*kernel[1]+tmp[6367]*kernel[2]+tmp[6465]*kernel[3]+tmp[6466]*kernel[4]+tmp[6467]*kernel[5]+tmp[6565]*kernel[6]+tmp[6566]*kernel[7]+tmp[6567]*kernel[8];
				ans[6467]<=tmp[6366]*kernel[0]+tmp[6367]*kernel[1]+tmp[6368]*kernel[2]+tmp[6466]*kernel[3]+tmp[6467]*kernel[4]+tmp[6468]*kernel[5]+tmp[6566]*kernel[6]+tmp[6567]*kernel[7]+tmp[6568]*kernel[8];
				ans[6468]<=tmp[6367]*kernel[0]+tmp[6368]*kernel[1]+tmp[6369]*kernel[2]+tmp[6467]*kernel[3]+tmp[6468]*kernel[4]+tmp[6469]*kernel[5]+tmp[6567]*kernel[6]+tmp[6568]*kernel[7]+tmp[6569]*kernel[8];
				ans[6469]<=tmp[6368]*kernel[0]+tmp[6369]*kernel[1]+tmp[6370]*kernel[2]+tmp[6468]*kernel[3]+tmp[6469]*kernel[4]+tmp[6470]*kernel[5]+tmp[6568]*kernel[6]+tmp[6569]*kernel[7]+tmp[6570]*kernel[8];
				ans[6470]<=tmp[6369]*kernel[0]+tmp[6370]*kernel[1]+tmp[6371]*kernel[2]+tmp[6469]*kernel[3]+tmp[6470]*kernel[4]+tmp[6471]*kernel[5]+tmp[6569]*kernel[6]+tmp[6570]*kernel[7]+tmp[6571]*kernel[8];
				ans[6471]<=tmp[6370]*kernel[0]+tmp[6371]*kernel[1]+tmp[6372]*kernel[2]+tmp[6470]*kernel[3]+tmp[6471]*kernel[4]+tmp[6472]*kernel[5]+tmp[6570]*kernel[6]+tmp[6571]*kernel[7]+tmp[6572]*kernel[8];
				ans[6472]<=tmp[6371]*kernel[0]+tmp[6372]*kernel[1]+tmp[6373]*kernel[2]+tmp[6471]*kernel[3]+tmp[6472]*kernel[4]+tmp[6473]*kernel[5]+tmp[6571]*kernel[6]+tmp[6572]*kernel[7]+tmp[6573]*kernel[8];
				ans[6473]<=tmp[6372]*kernel[0]+tmp[6373]*kernel[1]+tmp[6374]*kernel[2]+tmp[6472]*kernel[3]+tmp[6473]*kernel[4]+tmp[6474]*kernel[5]+tmp[6572]*kernel[6]+tmp[6573]*kernel[7]+tmp[6574]*kernel[8];
				ans[6474]<=tmp[6373]*kernel[0]+tmp[6374]*kernel[1]+tmp[6375]*kernel[2]+tmp[6473]*kernel[3]+tmp[6474]*kernel[4]+tmp[6475]*kernel[5]+tmp[6573]*kernel[6]+tmp[6574]*kernel[7]+tmp[6575]*kernel[8];
				ans[6475]<=tmp[6374]*kernel[0]+tmp[6375]*kernel[1]+tmp[6376]*kernel[2]+tmp[6474]*kernel[3]+tmp[6475]*kernel[4]+tmp[6476]*kernel[5]+tmp[6574]*kernel[6]+tmp[6575]*kernel[7]+tmp[6576]*kernel[8];
				ans[6476]<=tmp[6375]*kernel[0]+tmp[6376]*kernel[1]+tmp[6377]*kernel[2]+tmp[6475]*kernel[3]+tmp[6476]*kernel[4]+tmp[6477]*kernel[5]+tmp[6575]*kernel[6]+tmp[6576]*kernel[7]+tmp[6577]*kernel[8];
				ans[6477]<=tmp[6376]*kernel[0]+tmp[6377]*kernel[1]+tmp[6378]*kernel[2]+tmp[6476]*kernel[3]+tmp[6477]*kernel[4]+tmp[6478]*kernel[5]+tmp[6576]*kernel[6]+tmp[6577]*kernel[7]+tmp[6578]*kernel[8];
				ans[6478]<=tmp[6377]*kernel[0]+tmp[6378]*kernel[1]+tmp[6379]*kernel[2]+tmp[6477]*kernel[3]+tmp[6478]*kernel[4]+tmp[6479]*kernel[5]+tmp[6577]*kernel[6]+tmp[6578]*kernel[7]+tmp[6579]*kernel[8];
				ans[6479]<=tmp[6378]*kernel[0]+tmp[6379]*kernel[1]+tmp[6380]*kernel[2]+tmp[6478]*kernel[3]+tmp[6479]*kernel[4]+tmp[6480]*kernel[5]+tmp[6578]*kernel[6]+tmp[6579]*kernel[7]+tmp[6580]*kernel[8];
				ans[6480]<=tmp[6379]*kernel[0]+tmp[6380]*kernel[1]+tmp[6381]*kernel[2]+tmp[6479]*kernel[3]+tmp[6480]*kernel[4]+tmp[6481]*kernel[5]+tmp[6579]*kernel[6]+tmp[6580]*kernel[7]+tmp[6581]*kernel[8];
				ans[6481]<=tmp[6380]*kernel[0]+tmp[6381]*kernel[1]+tmp[6382]*kernel[2]+tmp[6480]*kernel[3]+tmp[6481]*kernel[4]+tmp[6482]*kernel[5]+tmp[6580]*kernel[6]+tmp[6581]*kernel[7]+tmp[6582]*kernel[8];
				ans[6482]<=tmp[6381]*kernel[0]+tmp[6382]*kernel[1]+tmp[6383]*kernel[2]+tmp[6481]*kernel[3]+tmp[6482]*kernel[4]+tmp[6483]*kernel[5]+tmp[6581]*kernel[6]+tmp[6582]*kernel[7]+tmp[6583]*kernel[8];
				ans[6483]<=tmp[6382]*kernel[0]+tmp[6383]*kernel[1]+tmp[6384]*kernel[2]+tmp[6482]*kernel[3]+tmp[6483]*kernel[4]+tmp[6484]*kernel[5]+tmp[6582]*kernel[6]+tmp[6583]*kernel[7]+tmp[6584]*kernel[8];
				ans[6484]<=tmp[6383]*kernel[0]+tmp[6384]*kernel[1]+tmp[6385]*kernel[2]+tmp[6483]*kernel[3]+tmp[6484]*kernel[4]+tmp[6485]*kernel[5]+tmp[6583]*kernel[6]+tmp[6584]*kernel[7]+tmp[6585]*kernel[8];
				ans[6485]<=tmp[6384]*kernel[0]+tmp[6385]*kernel[1]+tmp[6386]*kernel[2]+tmp[6484]*kernel[3]+tmp[6485]*kernel[4]+tmp[6486]*kernel[5]+tmp[6584]*kernel[6]+tmp[6585]*kernel[7]+tmp[6586]*kernel[8];
				ans[6486]<=tmp[6385]*kernel[0]+tmp[6386]*kernel[1]+tmp[6387]*kernel[2]+tmp[6485]*kernel[3]+tmp[6486]*kernel[4]+tmp[6487]*kernel[5]+tmp[6585]*kernel[6]+tmp[6586]*kernel[7]+tmp[6587]*kernel[8];
				ans[6487]<=tmp[6386]*kernel[0]+tmp[6387]*kernel[1]+tmp[6388]*kernel[2]+tmp[6486]*kernel[3]+tmp[6487]*kernel[4]+tmp[6488]*kernel[5]+tmp[6586]*kernel[6]+tmp[6587]*kernel[7]+tmp[6588]*kernel[8];
				ans[6488]<=tmp[6387]*kernel[0]+tmp[6388]*kernel[1]+tmp[6389]*kernel[2]+tmp[6487]*kernel[3]+tmp[6488]*kernel[4]+tmp[6489]*kernel[5]+tmp[6587]*kernel[6]+tmp[6588]*kernel[7]+tmp[6589]*kernel[8];
				ans[6489]<=tmp[6388]*kernel[0]+tmp[6389]*kernel[1]+tmp[6390]*kernel[2]+tmp[6488]*kernel[3]+tmp[6489]*kernel[4]+tmp[6490]*kernel[5]+tmp[6588]*kernel[6]+tmp[6589]*kernel[7]+tmp[6590]*kernel[8];
				ans[6490]<=tmp[6389]*kernel[0]+tmp[6390]*kernel[1]+tmp[6391]*kernel[2]+tmp[6489]*kernel[3]+tmp[6490]*kernel[4]+tmp[6491]*kernel[5]+tmp[6589]*kernel[6]+tmp[6590]*kernel[7]+tmp[6591]*kernel[8];
				ans[6491]<=tmp[6390]*kernel[0]+tmp[6391]*kernel[1]+tmp[6392]*kernel[2]+tmp[6490]*kernel[3]+tmp[6491]*kernel[4]+tmp[6492]*kernel[5]+tmp[6590]*kernel[6]+tmp[6591]*kernel[7]+tmp[6592]*kernel[8];
				ans[6492]<=tmp[6391]*kernel[0]+tmp[6392]*kernel[1]+tmp[6393]*kernel[2]+tmp[6491]*kernel[3]+tmp[6492]*kernel[4]+tmp[6493]*kernel[5]+tmp[6591]*kernel[6]+tmp[6592]*kernel[7]+tmp[6593]*kernel[8];
				ans[6493]<=tmp[6392]*kernel[0]+tmp[6393]*kernel[1]+tmp[6394]*kernel[2]+tmp[6492]*kernel[3]+tmp[6493]*kernel[4]+tmp[6494]*kernel[5]+tmp[6592]*kernel[6]+tmp[6593]*kernel[7]+tmp[6594]*kernel[8];
				ans[6494]<=tmp[6393]*kernel[0]+tmp[6394]*kernel[1]+tmp[6395]*kernel[2]+tmp[6493]*kernel[3]+tmp[6494]*kernel[4]+tmp[6495]*kernel[5]+tmp[6593]*kernel[6]+tmp[6594]*kernel[7]+tmp[6595]*kernel[8];
				ans[6495]<=tmp[6394]*kernel[0]+tmp[6395]*kernel[1]+tmp[6396]*kernel[2]+tmp[6494]*kernel[3]+tmp[6495]*kernel[4]+tmp[6496]*kernel[5]+tmp[6594]*kernel[6]+tmp[6595]*kernel[7]+tmp[6596]*kernel[8];
				ans[6496]<=tmp[6395]*kernel[0]+tmp[6396]*kernel[1]+tmp[6397]*kernel[2]+tmp[6495]*kernel[3]+tmp[6496]*kernel[4]+tmp[6497]*kernel[5]+tmp[6595]*kernel[6]+tmp[6596]*kernel[7]+tmp[6597]*kernel[8];
				ans[6497]<=tmp[6396]*kernel[0]+tmp[6397]*kernel[1]+tmp[6398]*kernel[2]+tmp[6496]*kernel[3]+tmp[6497]*kernel[4]+tmp[6498]*kernel[5]+tmp[6596]*kernel[6]+tmp[6597]*kernel[7]+tmp[6598]*kernel[8];
				ans[6498]<=tmp[6397]*kernel[0]+tmp[6398]*kernel[1]+tmp[6399]*kernel[2]+tmp[6497]*kernel[3]+tmp[6498]*kernel[4]+tmp[6499]*kernel[5]+tmp[6597]*kernel[6]+tmp[6598]*kernel[7]+tmp[6599]*kernel[8];
				ans[6499]<=tmp[6398]*kernel[0]+tmp[6399]*kernel[1]+tmp[6498]*kernel[3]+tmp[6499]*kernel[4]+tmp[6598]*kernel[6]+tmp[6599]*kernel[7];
				ans[6500]<=tmp[6400]*kernel[1]+tmp[6401]*kernel[2]+tmp[6500]*kernel[4]+tmp[6501]*kernel[5]+tmp[6600]*kernel[7]+tmp[6601]*kernel[8];
				ans[6501]<=tmp[6400]*kernel[0]+tmp[6401]*kernel[1]+tmp[6402]*kernel[2]+tmp[6500]*kernel[3]+tmp[6501]*kernel[4]+tmp[6502]*kernel[5]+tmp[6600]*kernel[6]+tmp[6601]*kernel[7]+tmp[6602]*kernel[8];
				ans[6502]<=tmp[6401]*kernel[0]+tmp[6402]*kernel[1]+tmp[6403]*kernel[2]+tmp[6501]*kernel[3]+tmp[6502]*kernel[4]+tmp[6503]*kernel[5]+tmp[6601]*kernel[6]+tmp[6602]*kernel[7]+tmp[6603]*kernel[8];
				ans[6503]<=tmp[6402]*kernel[0]+tmp[6403]*kernel[1]+tmp[6404]*kernel[2]+tmp[6502]*kernel[3]+tmp[6503]*kernel[4]+tmp[6504]*kernel[5]+tmp[6602]*kernel[6]+tmp[6603]*kernel[7]+tmp[6604]*kernel[8];
				ans[6504]<=tmp[6403]*kernel[0]+tmp[6404]*kernel[1]+tmp[6405]*kernel[2]+tmp[6503]*kernel[3]+tmp[6504]*kernel[4]+tmp[6505]*kernel[5]+tmp[6603]*kernel[6]+tmp[6604]*kernel[7]+tmp[6605]*kernel[8];
				ans[6505]<=tmp[6404]*kernel[0]+tmp[6405]*kernel[1]+tmp[6406]*kernel[2]+tmp[6504]*kernel[3]+tmp[6505]*kernel[4]+tmp[6506]*kernel[5]+tmp[6604]*kernel[6]+tmp[6605]*kernel[7]+tmp[6606]*kernel[8];
				ans[6506]<=tmp[6405]*kernel[0]+tmp[6406]*kernel[1]+tmp[6407]*kernel[2]+tmp[6505]*kernel[3]+tmp[6506]*kernel[4]+tmp[6507]*kernel[5]+tmp[6605]*kernel[6]+tmp[6606]*kernel[7]+tmp[6607]*kernel[8];
				ans[6507]<=tmp[6406]*kernel[0]+tmp[6407]*kernel[1]+tmp[6408]*kernel[2]+tmp[6506]*kernel[3]+tmp[6507]*kernel[4]+tmp[6508]*kernel[5]+tmp[6606]*kernel[6]+tmp[6607]*kernel[7]+tmp[6608]*kernel[8];
				ans[6508]<=tmp[6407]*kernel[0]+tmp[6408]*kernel[1]+tmp[6409]*kernel[2]+tmp[6507]*kernel[3]+tmp[6508]*kernel[4]+tmp[6509]*kernel[5]+tmp[6607]*kernel[6]+tmp[6608]*kernel[7]+tmp[6609]*kernel[8];
				ans[6509]<=tmp[6408]*kernel[0]+tmp[6409]*kernel[1]+tmp[6410]*kernel[2]+tmp[6508]*kernel[3]+tmp[6509]*kernel[4]+tmp[6510]*kernel[5]+tmp[6608]*kernel[6]+tmp[6609]*kernel[7]+tmp[6610]*kernel[8];
				ans[6510]<=tmp[6409]*kernel[0]+tmp[6410]*kernel[1]+tmp[6411]*kernel[2]+tmp[6509]*kernel[3]+tmp[6510]*kernel[4]+tmp[6511]*kernel[5]+tmp[6609]*kernel[6]+tmp[6610]*kernel[7]+tmp[6611]*kernel[8];
				ans[6511]<=tmp[6410]*kernel[0]+tmp[6411]*kernel[1]+tmp[6412]*kernel[2]+tmp[6510]*kernel[3]+tmp[6511]*kernel[4]+tmp[6512]*kernel[5]+tmp[6610]*kernel[6]+tmp[6611]*kernel[7]+tmp[6612]*kernel[8];
				ans[6512]<=tmp[6411]*kernel[0]+tmp[6412]*kernel[1]+tmp[6413]*kernel[2]+tmp[6511]*kernel[3]+tmp[6512]*kernel[4]+tmp[6513]*kernel[5]+tmp[6611]*kernel[6]+tmp[6612]*kernel[7]+tmp[6613]*kernel[8];
				ans[6513]<=tmp[6412]*kernel[0]+tmp[6413]*kernel[1]+tmp[6414]*kernel[2]+tmp[6512]*kernel[3]+tmp[6513]*kernel[4]+tmp[6514]*kernel[5]+tmp[6612]*kernel[6]+tmp[6613]*kernel[7]+tmp[6614]*kernel[8];
				ans[6514]<=tmp[6413]*kernel[0]+tmp[6414]*kernel[1]+tmp[6415]*kernel[2]+tmp[6513]*kernel[3]+tmp[6514]*kernel[4]+tmp[6515]*kernel[5]+tmp[6613]*kernel[6]+tmp[6614]*kernel[7]+tmp[6615]*kernel[8];
				ans[6515]<=tmp[6414]*kernel[0]+tmp[6415]*kernel[1]+tmp[6416]*kernel[2]+tmp[6514]*kernel[3]+tmp[6515]*kernel[4]+tmp[6516]*kernel[5]+tmp[6614]*kernel[6]+tmp[6615]*kernel[7]+tmp[6616]*kernel[8];
				ans[6516]<=tmp[6415]*kernel[0]+tmp[6416]*kernel[1]+tmp[6417]*kernel[2]+tmp[6515]*kernel[3]+tmp[6516]*kernel[4]+tmp[6517]*kernel[5]+tmp[6615]*kernel[6]+tmp[6616]*kernel[7]+tmp[6617]*kernel[8];
				ans[6517]<=tmp[6416]*kernel[0]+tmp[6417]*kernel[1]+tmp[6418]*kernel[2]+tmp[6516]*kernel[3]+tmp[6517]*kernel[4]+tmp[6518]*kernel[5]+tmp[6616]*kernel[6]+tmp[6617]*kernel[7]+tmp[6618]*kernel[8];
				ans[6518]<=tmp[6417]*kernel[0]+tmp[6418]*kernel[1]+tmp[6419]*kernel[2]+tmp[6517]*kernel[3]+tmp[6518]*kernel[4]+tmp[6519]*kernel[5]+tmp[6617]*kernel[6]+tmp[6618]*kernel[7]+tmp[6619]*kernel[8];
				ans[6519]<=tmp[6418]*kernel[0]+tmp[6419]*kernel[1]+tmp[6420]*kernel[2]+tmp[6518]*kernel[3]+tmp[6519]*kernel[4]+tmp[6520]*kernel[5]+tmp[6618]*kernel[6]+tmp[6619]*kernel[7]+tmp[6620]*kernel[8];
				ans[6520]<=tmp[6419]*kernel[0]+tmp[6420]*kernel[1]+tmp[6421]*kernel[2]+tmp[6519]*kernel[3]+tmp[6520]*kernel[4]+tmp[6521]*kernel[5]+tmp[6619]*kernel[6]+tmp[6620]*kernel[7]+tmp[6621]*kernel[8];
				ans[6521]<=tmp[6420]*kernel[0]+tmp[6421]*kernel[1]+tmp[6422]*kernel[2]+tmp[6520]*kernel[3]+tmp[6521]*kernel[4]+tmp[6522]*kernel[5]+tmp[6620]*kernel[6]+tmp[6621]*kernel[7]+tmp[6622]*kernel[8];
				ans[6522]<=tmp[6421]*kernel[0]+tmp[6422]*kernel[1]+tmp[6423]*kernel[2]+tmp[6521]*kernel[3]+tmp[6522]*kernel[4]+tmp[6523]*kernel[5]+tmp[6621]*kernel[6]+tmp[6622]*kernel[7]+tmp[6623]*kernel[8];
				ans[6523]<=tmp[6422]*kernel[0]+tmp[6423]*kernel[1]+tmp[6424]*kernel[2]+tmp[6522]*kernel[3]+tmp[6523]*kernel[4]+tmp[6524]*kernel[5]+tmp[6622]*kernel[6]+tmp[6623]*kernel[7]+tmp[6624]*kernel[8];
				ans[6524]<=tmp[6423]*kernel[0]+tmp[6424]*kernel[1]+tmp[6425]*kernel[2]+tmp[6523]*kernel[3]+tmp[6524]*kernel[4]+tmp[6525]*kernel[5]+tmp[6623]*kernel[6]+tmp[6624]*kernel[7]+tmp[6625]*kernel[8];
				ans[6525]<=tmp[6424]*kernel[0]+tmp[6425]*kernel[1]+tmp[6426]*kernel[2]+tmp[6524]*kernel[3]+tmp[6525]*kernel[4]+tmp[6526]*kernel[5]+tmp[6624]*kernel[6]+tmp[6625]*kernel[7]+tmp[6626]*kernel[8];
				ans[6526]<=tmp[6425]*kernel[0]+tmp[6426]*kernel[1]+tmp[6427]*kernel[2]+tmp[6525]*kernel[3]+tmp[6526]*kernel[4]+tmp[6527]*kernel[5]+tmp[6625]*kernel[6]+tmp[6626]*kernel[7]+tmp[6627]*kernel[8];
				ans[6527]<=tmp[6426]*kernel[0]+tmp[6427]*kernel[1]+tmp[6428]*kernel[2]+tmp[6526]*kernel[3]+tmp[6527]*kernel[4]+tmp[6528]*kernel[5]+tmp[6626]*kernel[6]+tmp[6627]*kernel[7]+tmp[6628]*kernel[8];
				ans[6528]<=tmp[6427]*kernel[0]+tmp[6428]*kernel[1]+tmp[6429]*kernel[2]+tmp[6527]*kernel[3]+tmp[6528]*kernel[4]+tmp[6529]*kernel[5]+tmp[6627]*kernel[6]+tmp[6628]*kernel[7]+tmp[6629]*kernel[8];
				ans[6529]<=tmp[6428]*kernel[0]+tmp[6429]*kernel[1]+tmp[6430]*kernel[2]+tmp[6528]*kernel[3]+tmp[6529]*kernel[4]+tmp[6530]*kernel[5]+tmp[6628]*kernel[6]+tmp[6629]*kernel[7]+tmp[6630]*kernel[8];
				ans[6530]<=tmp[6429]*kernel[0]+tmp[6430]*kernel[1]+tmp[6431]*kernel[2]+tmp[6529]*kernel[3]+tmp[6530]*kernel[4]+tmp[6531]*kernel[5]+tmp[6629]*kernel[6]+tmp[6630]*kernel[7]+tmp[6631]*kernel[8];
				ans[6531]<=tmp[6430]*kernel[0]+tmp[6431]*kernel[1]+tmp[6432]*kernel[2]+tmp[6530]*kernel[3]+tmp[6531]*kernel[4]+tmp[6532]*kernel[5]+tmp[6630]*kernel[6]+tmp[6631]*kernel[7]+tmp[6632]*kernel[8];
				ans[6532]<=tmp[6431]*kernel[0]+tmp[6432]*kernel[1]+tmp[6433]*kernel[2]+tmp[6531]*kernel[3]+tmp[6532]*kernel[4]+tmp[6533]*kernel[5]+tmp[6631]*kernel[6]+tmp[6632]*kernel[7]+tmp[6633]*kernel[8];
				ans[6533]<=tmp[6432]*kernel[0]+tmp[6433]*kernel[1]+tmp[6434]*kernel[2]+tmp[6532]*kernel[3]+tmp[6533]*kernel[4]+tmp[6534]*kernel[5]+tmp[6632]*kernel[6]+tmp[6633]*kernel[7]+tmp[6634]*kernel[8];
				ans[6534]<=tmp[6433]*kernel[0]+tmp[6434]*kernel[1]+tmp[6435]*kernel[2]+tmp[6533]*kernel[3]+tmp[6534]*kernel[4]+tmp[6535]*kernel[5]+tmp[6633]*kernel[6]+tmp[6634]*kernel[7]+tmp[6635]*kernel[8];
				ans[6535]<=tmp[6434]*kernel[0]+tmp[6435]*kernel[1]+tmp[6436]*kernel[2]+tmp[6534]*kernel[3]+tmp[6535]*kernel[4]+tmp[6536]*kernel[5]+tmp[6634]*kernel[6]+tmp[6635]*kernel[7]+tmp[6636]*kernel[8];
				ans[6536]<=tmp[6435]*kernel[0]+tmp[6436]*kernel[1]+tmp[6437]*kernel[2]+tmp[6535]*kernel[3]+tmp[6536]*kernel[4]+tmp[6537]*kernel[5]+tmp[6635]*kernel[6]+tmp[6636]*kernel[7]+tmp[6637]*kernel[8];
				ans[6537]<=tmp[6436]*kernel[0]+tmp[6437]*kernel[1]+tmp[6438]*kernel[2]+tmp[6536]*kernel[3]+tmp[6537]*kernel[4]+tmp[6538]*kernel[5]+tmp[6636]*kernel[6]+tmp[6637]*kernel[7]+tmp[6638]*kernel[8];
				ans[6538]<=tmp[6437]*kernel[0]+tmp[6438]*kernel[1]+tmp[6439]*kernel[2]+tmp[6537]*kernel[3]+tmp[6538]*kernel[4]+tmp[6539]*kernel[5]+tmp[6637]*kernel[6]+tmp[6638]*kernel[7]+tmp[6639]*kernel[8];
				ans[6539]<=tmp[6438]*kernel[0]+tmp[6439]*kernel[1]+tmp[6440]*kernel[2]+tmp[6538]*kernel[3]+tmp[6539]*kernel[4]+tmp[6540]*kernel[5]+tmp[6638]*kernel[6]+tmp[6639]*kernel[7]+tmp[6640]*kernel[8];
				ans[6540]<=tmp[6439]*kernel[0]+tmp[6440]*kernel[1]+tmp[6441]*kernel[2]+tmp[6539]*kernel[3]+tmp[6540]*kernel[4]+tmp[6541]*kernel[5]+tmp[6639]*kernel[6]+tmp[6640]*kernel[7]+tmp[6641]*kernel[8];
				ans[6541]<=tmp[6440]*kernel[0]+tmp[6441]*kernel[1]+tmp[6442]*kernel[2]+tmp[6540]*kernel[3]+tmp[6541]*kernel[4]+tmp[6542]*kernel[5]+tmp[6640]*kernel[6]+tmp[6641]*kernel[7]+tmp[6642]*kernel[8];
				ans[6542]<=tmp[6441]*kernel[0]+tmp[6442]*kernel[1]+tmp[6443]*kernel[2]+tmp[6541]*kernel[3]+tmp[6542]*kernel[4]+tmp[6543]*kernel[5]+tmp[6641]*kernel[6]+tmp[6642]*kernel[7]+tmp[6643]*kernel[8];
				ans[6543]<=tmp[6442]*kernel[0]+tmp[6443]*kernel[1]+tmp[6444]*kernel[2]+tmp[6542]*kernel[3]+tmp[6543]*kernel[4]+tmp[6544]*kernel[5]+tmp[6642]*kernel[6]+tmp[6643]*kernel[7]+tmp[6644]*kernel[8];
				ans[6544]<=tmp[6443]*kernel[0]+tmp[6444]*kernel[1]+tmp[6445]*kernel[2]+tmp[6543]*kernel[3]+tmp[6544]*kernel[4]+tmp[6545]*kernel[5]+tmp[6643]*kernel[6]+tmp[6644]*kernel[7]+tmp[6645]*kernel[8];
				ans[6545]<=tmp[6444]*kernel[0]+tmp[6445]*kernel[1]+tmp[6446]*kernel[2]+tmp[6544]*kernel[3]+tmp[6545]*kernel[4]+tmp[6546]*kernel[5]+tmp[6644]*kernel[6]+tmp[6645]*kernel[7]+tmp[6646]*kernel[8];
				ans[6546]<=tmp[6445]*kernel[0]+tmp[6446]*kernel[1]+tmp[6447]*kernel[2]+tmp[6545]*kernel[3]+tmp[6546]*kernel[4]+tmp[6547]*kernel[5]+tmp[6645]*kernel[6]+tmp[6646]*kernel[7]+tmp[6647]*kernel[8];
				ans[6547]<=tmp[6446]*kernel[0]+tmp[6447]*kernel[1]+tmp[6448]*kernel[2]+tmp[6546]*kernel[3]+tmp[6547]*kernel[4]+tmp[6548]*kernel[5]+tmp[6646]*kernel[6]+tmp[6647]*kernel[7]+tmp[6648]*kernel[8];
				ans[6548]<=tmp[6447]*kernel[0]+tmp[6448]*kernel[1]+tmp[6449]*kernel[2]+tmp[6547]*kernel[3]+tmp[6548]*kernel[4]+tmp[6549]*kernel[5]+tmp[6647]*kernel[6]+tmp[6648]*kernel[7]+tmp[6649]*kernel[8];
				ans[6549]<=tmp[6448]*kernel[0]+tmp[6449]*kernel[1]+tmp[6450]*kernel[2]+tmp[6548]*kernel[3]+tmp[6549]*kernel[4]+tmp[6550]*kernel[5]+tmp[6648]*kernel[6]+tmp[6649]*kernel[7]+tmp[6650]*kernel[8];
				ans[6550]<=tmp[6449]*kernel[0]+tmp[6450]*kernel[1]+tmp[6451]*kernel[2]+tmp[6549]*kernel[3]+tmp[6550]*kernel[4]+tmp[6551]*kernel[5]+tmp[6649]*kernel[6]+tmp[6650]*kernel[7]+tmp[6651]*kernel[8];
				ans[6551]<=tmp[6450]*kernel[0]+tmp[6451]*kernel[1]+tmp[6452]*kernel[2]+tmp[6550]*kernel[3]+tmp[6551]*kernel[4]+tmp[6552]*kernel[5]+tmp[6650]*kernel[6]+tmp[6651]*kernel[7]+tmp[6652]*kernel[8];
				ans[6552]<=tmp[6451]*kernel[0]+tmp[6452]*kernel[1]+tmp[6453]*kernel[2]+tmp[6551]*kernel[3]+tmp[6552]*kernel[4]+tmp[6553]*kernel[5]+tmp[6651]*kernel[6]+tmp[6652]*kernel[7]+tmp[6653]*kernel[8];
				ans[6553]<=tmp[6452]*kernel[0]+tmp[6453]*kernel[1]+tmp[6454]*kernel[2]+tmp[6552]*kernel[3]+tmp[6553]*kernel[4]+tmp[6554]*kernel[5]+tmp[6652]*kernel[6]+tmp[6653]*kernel[7]+tmp[6654]*kernel[8];
				ans[6554]<=tmp[6453]*kernel[0]+tmp[6454]*kernel[1]+tmp[6455]*kernel[2]+tmp[6553]*kernel[3]+tmp[6554]*kernel[4]+tmp[6555]*kernel[5]+tmp[6653]*kernel[6]+tmp[6654]*kernel[7]+tmp[6655]*kernel[8];
				ans[6555]<=tmp[6454]*kernel[0]+tmp[6455]*kernel[1]+tmp[6456]*kernel[2]+tmp[6554]*kernel[3]+tmp[6555]*kernel[4]+tmp[6556]*kernel[5]+tmp[6654]*kernel[6]+tmp[6655]*kernel[7]+tmp[6656]*kernel[8];
				ans[6556]<=tmp[6455]*kernel[0]+tmp[6456]*kernel[1]+tmp[6457]*kernel[2]+tmp[6555]*kernel[3]+tmp[6556]*kernel[4]+tmp[6557]*kernel[5]+tmp[6655]*kernel[6]+tmp[6656]*kernel[7]+tmp[6657]*kernel[8];
				ans[6557]<=tmp[6456]*kernel[0]+tmp[6457]*kernel[1]+tmp[6458]*kernel[2]+tmp[6556]*kernel[3]+tmp[6557]*kernel[4]+tmp[6558]*kernel[5]+tmp[6656]*kernel[6]+tmp[6657]*kernel[7]+tmp[6658]*kernel[8];
				ans[6558]<=tmp[6457]*kernel[0]+tmp[6458]*kernel[1]+tmp[6459]*kernel[2]+tmp[6557]*kernel[3]+tmp[6558]*kernel[4]+tmp[6559]*kernel[5]+tmp[6657]*kernel[6]+tmp[6658]*kernel[7]+tmp[6659]*kernel[8];
				ans[6559]<=tmp[6458]*kernel[0]+tmp[6459]*kernel[1]+tmp[6460]*kernel[2]+tmp[6558]*kernel[3]+tmp[6559]*kernel[4]+tmp[6560]*kernel[5]+tmp[6658]*kernel[6]+tmp[6659]*kernel[7]+tmp[6660]*kernel[8];
				ans[6560]<=tmp[6459]*kernel[0]+tmp[6460]*kernel[1]+tmp[6461]*kernel[2]+tmp[6559]*kernel[3]+tmp[6560]*kernel[4]+tmp[6561]*kernel[5]+tmp[6659]*kernel[6]+tmp[6660]*kernel[7]+tmp[6661]*kernel[8];
				ans[6561]<=tmp[6460]*kernel[0]+tmp[6461]*kernel[1]+tmp[6462]*kernel[2]+tmp[6560]*kernel[3]+tmp[6561]*kernel[4]+tmp[6562]*kernel[5]+tmp[6660]*kernel[6]+tmp[6661]*kernel[7]+tmp[6662]*kernel[8];
				ans[6562]<=tmp[6461]*kernel[0]+tmp[6462]*kernel[1]+tmp[6463]*kernel[2]+tmp[6561]*kernel[3]+tmp[6562]*kernel[4]+tmp[6563]*kernel[5]+tmp[6661]*kernel[6]+tmp[6662]*kernel[7]+tmp[6663]*kernel[8];
				ans[6563]<=tmp[6462]*kernel[0]+tmp[6463]*kernel[1]+tmp[6464]*kernel[2]+tmp[6562]*kernel[3]+tmp[6563]*kernel[4]+tmp[6564]*kernel[5]+tmp[6662]*kernel[6]+tmp[6663]*kernel[7]+tmp[6664]*kernel[8];
				ans[6564]<=tmp[6463]*kernel[0]+tmp[6464]*kernel[1]+tmp[6465]*kernel[2]+tmp[6563]*kernel[3]+tmp[6564]*kernel[4]+tmp[6565]*kernel[5]+tmp[6663]*kernel[6]+tmp[6664]*kernel[7]+tmp[6665]*kernel[8];
				ans[6565]<=tmp[6464]*kernel[0]+tmp[6465]*kernel[1]+tmp[6466]*kernel[2]+tmp[6564]*kernel[3]+tmp[6565]*kernel[4]+tmp[6566]*kernel[5]+tmp[6664]*kernel[6]+tmp[6665]*kernel[7]+tmp[6666]*kernel[8];
				ans[6566]<=tmp[6465]*kernel[0]+tmp[6466]*kernel[1]+tmp[6467]*kernel[2]+tmp[6565]*kernel[3]+tmp[6566]*kernel[4]+tmp[6567]*kernel[5]+tmp[6665]*kernel[6]+tmp[6666]*kernel[7]+tmp[6667]*kernel[8];
				ans[6567]<=tmp[6466]*kernel[0]+tmp[6467]*kernel[1]+tmp[6468]*kernel[2]+tmp[6566]*kernel[3]+tmp[6567]*kernel[4]+tmp[6568]*kernel[5]+tmp[6666]*kernel[6]+tmp[6667]*kernel[7]+tmp[6668]*kernel[8];
				ans[6568]<=tmp[6467]*kernel[0]+tmp[6468]*kernel[1]+tmp[6469]*kernel[2]+tmp[6567]*kernel[3]+tmp[6568]*kernel[4]+tmp[6569]*kernel[5]+tmp[6667]*kernel[6]+tmp[6668]*kernel[7]+tmp[6669]*kernel[8];
				ans[6569]<=tmp[6468]*kernel[0]+tmp[6469]*kernel[1]+tmp[6470]*kernel[2]+tmp[6568]*kernel[3]+tmp[6569]*kernel[4]+tmp[6570]*kernel[5]+tmp[6668]*kernel[6]+tmp[6669]*kernel[7]+tmp[6670]*kernel[8];
				ans[6570]<=tmp[6469]*kernel[0]+tmp[6470]*kernel[1]+tmp[6471]*kernel[2]+tmp[6569]*kernel[3]+tmp[6570]*kernel[4]+tmp[6571]*kernel[5]+tmp[6669]*kernel[6]+tmp[6670]*kernel[7]+tmp[6671]*kernel[8];
				ans[6571]<=tmp[6470]*kernel[0]+tmp[6471]*kernel[1]+tmp[6472]*kernel[2]+tmp[6570]*kernel[3]+tmp[6571]*kernel[4]+tmp[6572]*kernel[5]+tmp[6670]*kernel[6]+tmp[6671]*kernel[7]+tmp[6672]*kernel[8];
				ans[6572]<=tmp[6471]*kernel[0]+tmp[6472]*kernel[1]+tmp[6473]*kernel[2]+tmp[6571]*kernel[3]+tmp[6572]*kernel[4]+tmp[6573]*kernel[5]+tmp[6671]*kernel[6]+tmp[6672]*kernel[7]+tmp[6673]*kernel[8];
				ans[6573]<=tmp[6472]*kernel[0]+tmp[6473]*kernel[1]+tmp[6474]*kernel[2]+tmp[6572]*kernel[3]+tmp[6573]*kernel[4]+tmp[6574]*kernel[5]+tmp[6672]*kernel[6]+tmp[6673]*kernel[7]+tmp[6674]*kernel[8];
				ans[6574]<=tmp[6473]*kernel[0]+tmp[6474]*kernel[1]+tmp[6475]*kernel[2]+tmp[6573]*kernel[3]+tmp[6574]*kernel[4]+tmp[6575]*kernel[5]+tmp[6673]*kernel[6]+tmp[6674]*kernel[7]+tmp[6675]*kernel[8];
				ans[6575]<=tmp[6474]*kernel[0]+tmp[6475]*kernel[1]+tmp[6476]*kernel[2]+tmp[6574]*kernel[3]+tmp[6575]*kernel[4]+tmp[6576]*kernel[5]+tmp[6674]*kernel[6]+tmp[6675]*kernel[7]+tmp[6676]*kernel[8];
				ans[6576]<=tmp[6475]*kernel[0]+tmp[6476]*kernel[1]+tmp[6477]*kernel[2]+tmp[6575]*kernel[3]+tmp[6576]*kernel[4]+tmp[6577]*kernel[5]+tmp[6675]*kernel[6]+tmp[6676]*kernel[7]+tmp[6677]*kernel[8];
				ans[6577]<=tmp[6476]*kernel[0]+tmp[6477]*kernel[1]+tmp[6478]*kernel[2]+tmp[6576]*kernel[3]+tmp[6577]*kernel[4]+tmp[6578]*kernel[5]+tmp[6676]*kernel[6]+tmp[6677]*kernel[7]+tmp[6678]*kernel[8];
				ans[6578]<=tmp[6477]*kernel[0]+tmp[6478]*kernel[1]+tmp[6479]*kernel[2]+tmp[6577]*kernel[3]+tmp[6578]*kernel[4]+tmp[6579]*kernel[5]+tmp[6677]*kernel[6]+tmp[6678]*kernel[7]+tmp[6679]*kernel[8];
				ans[6579]<=tmp[6478]*kernel[0]+tmp[6479]*kernel[1]+tmp[6480]*kernel[2]+tmp[6578]*kernel[3]+tmp[6579]*kernel[4]+tmp[6580]*kernel[5]+tmp[6678]*kernel[6]+tmp[6679]*kernel[7]+tmp[6680]*kernel[8];
				ans[6580]<=tmp[6479]*kernel[0]+tmp[6480]*kernel[1]+tmp[6481]*kernel[2]+tmp[6579]*kernel[3]+tmp[6580]*kernel[4]+tmp[6581]*kernel[5]+tmp[6679]*kernel[6]+tmp[6680]*kernel[7]+tmp[6681]*kernel[8];
				ans[6581]<=tmp[6480]*kernel[0]+tmp[6481]*kernel[1]+tmp[6482]*kernel[2]+tmp[6580]*kernel[3]+tmp[6581]*kernel[4]+tmp[6582]*kernel[5]+tmp[6680]*kernel[6]+tmp[6681]*kernel[7]+tmp[6682]*kernel[8];
				ans[6582]<=tmp[6481]*kernel[0]+tmp[6482]*kernel[1]+tmp[6483]*kernel[2]+tmp[6581]*kernel[3]+tmp[6582]*kernel[4]+tmp[6583]*kernel[5]+tmp[6681]*kernel[6]+tmp[6682]*kernel[7]+tmp[6683]*kernel[8];
				ans[6583]<=tmp[6482]*kernel[0]+tmp[6483]*kernel[1]+tmp[6484]*kernel[2]+tmp[6582]*kernel[3]+tmp[6583]*kernel[4]+tmp[6584]*kernel[5]+tmp[6682]*kernel[6]+tmp[6683]*kernel[7]+tmp[6684]*kernel[8];
				ans[6584]<=tmp[6483]*kernel[0]+tmp[6484]*kernel[1]+tmp[6485]*kernel[2]+tmp[6583]*kernel[3]+tmp[6584]*kernel[4]+tmp[6585]*kernel[5]+tmp[6683]*kernel[6]+tmp[6684]*kernel[7]+tmp[6685]*kernel[8];
				ans[6585]<=tmp[6484]*kernel[0]+tmp[6485]*kernel[1]+tmp[6486]*kernel[2]+tmp[6584]*kernel[3]+tmp[6585]*kernel[4]+tmp[6586]*kernel[5]+tmp[6684]*kernel[6]+tmp[6685]*kernel[7]+tmp[6686]*kernel[8];
				ans[6586]<=tmp[6485]*kernel[0]+tmp[6486]*kernel[1]+tmp[6487]*kernel[2]+tmp[6585]*kernel[3]+tmp[6586]*kernel[4]+tmp[6587]*kernel[5]+tmp[6685]*kernel[6]+tmp[6686]*kernel[7]+tmp[6687]*kernel[8];
				ans[6587]<=tmp[6486]*kernel[0]+tmp[6487]*kernel[1]+tmp[6488]*kernel[2]+tmp[6586]*kernel[3]+tmp[6587]*kernel[4]+tmp[6588]*kernel[5]+tmp[6686]*kernel[6]+tmp[6687]*kernel[7]+tmp[6688]*kernel[8];
				ans[6588]<=tmp[6487]*kernel[0]+tmp[6488]*kernel[1]+tmp[6489]*kernel[2]+tmp[6587]*kernel[3]+tmp[6588]*kernel[4]+tmp[6589]*kernel[5]+tmp[6687]*kernel[6]+tmp[6688]*kernel[7]+tmp[6689]*kernel[8];
				ans[6589]<=tmp[6488]*kernel[0]+tmp[6489]*kernel[1]+tmp[6490]*kernel[2]+tmp[6588]*kernel[3]+tmp[6589]*kernel[4]+tmp[6590]*kernel[5]+tmp[6688]*kernel[6]+tmp[6689]*kernel[7]+tmp[6690]*kernel[8];
				ans[6590]<=tmp[6489]*kernel[0]+tmp[6490]*kernel[1]+tmp[6491]*kernel[2]+tmp[6589]*kernel[3]+tmp[6590]*kernel[4]+tmp[6591]*kernel[5]+tmp[6689]*kernel[6]+tmp[6690]*kernel[7]+tmp[6691]*kernel[8];
				ans[6591]<=tmp[6490]*kernel[0]+tmp[6491]*kernel[1]+tmp[6492]*kernel[2]+tmp[6590]*kernel[3]+tmp[6591]*kernel[4]+tmp[6592]*kernel[5]+tmp[6690]*kernel[6]+tmp[6691]*kernel[7]+tmp[6692]*kernel[8];
				ans[6592]<=tmp[6491]*kernel[0]+tmp[6492]*kernel[1]+tmp[6493]*kernel[2]+tmp[6591]*kernel[3]+tmp[6592]*kernel[4]+tmp[6593]*kernel[5]+tmp[6691]*kernel[6]+tmp[6692]*kernel[7]+tmp[6693]*kernel[8];
				ans[6593]<=tmp[6492]*kernel[0]+tmp[6493]*kernel[1]+tmp[6494]*kernel[2]+tmp[6592]*kernel[3]+tmp[6593]*kernel[4]+tmp[6594]*kernel[5]+tmp[6692]*kernel[6]+tmp[6693]*kernel[7]+tmp[6694]*kernel[8];
				ans[6594]<=tmp[6493]*kernel[0]+tmp[6494]*kernel[1]+tmp[6495]*kernel[2]+tmp[6593]*kernel[3]+tmp[6594]*kernel[4]+tmp[6595]*kernel[5]+tmp[6693]*kernel[6]+tmp[6694]*kernel[7]+tmp[6695]*kernel[8];
				ans[6595]<=tmp[6494]*kernel[0]+tmp[6495]*kernel[1]+tmp[6496]*kernel[2]+tmp[6594]*kernel[3]+tmp[6595]*kernel[4]+tmp[6596]*kernel[5]+tmp[6694]*kernel[6]+tmp[6695]*kernel[7]+tmp[6696]*kernel[8];
				ans[6596]<=tmp[6495]*kernel[0]+tmp[6496]*kernel[1]+tmp[6497]*kernel[2]+tmp[6595]*kernel[3]+tmp[6596]*kernel[4]+tmp[6597]*kernel[5]+tmp[6695]*kernel[6]+tmp[6696]*kernel[7]+tmp[6697]*kernel[8];
				ans[6597]<=tmp[6496]*kernel[0]+tmp[6497]*kernel[1]+tmp[6498]*kernel[2]+tmp[6596]*kernel[3]+tmp[6597]*kernel[4]+tmp[6598]*kernel[5]+tmp[6696]*kernel[6]+tmp[6697]*kernel[7]+tmp[6698]*kernel[8];
				ans[6598]<=tmp[6497]*kernel[0]+tmp[6498]*kernel[1]+tmp[6499]*kernel[2]+tmp[6597]*kernel[3]+tmp[6598]*kernel[4]+tmp[6599]*kernel[5]+tmp[6697]*kernel[6]+tmp[6698]*kernel[7]+tmp[6699]*kernel[8];
				ans[6599]<=tmp[6498]*kernel[0]+tmp[6499]*kernel[1]+tmp[6598]*kernel[3]+tmp[6599]*kernel[4]+tmp[6698]*kernel[6]+tmp[6699]*kernel[7];
				ans[6600]<=tmp[6500]*kernel[1]+tmp[6501]*kernel[2]+tmp[6600]*kernel[4]+tmp[6601]*kernel[5]+tmp[6700]*kernel[7]+tmp[6701]*kernel[8];
				ans[6601]<=tmp[6500]*kernel[0]+tmp[6501]*kernel[1]+tmp[6502]*kernel[2]+tmp[6600]*kernel[3]+tmp[6601]*kernel[4]+tmp[6602]*kernel[5]+tmp[6700]*kernel[6]+tmp[6701]*kernel[7]+tmp[6702]*kernel[8];
				ans[6602]<=tmp[6501]*kernel[0]+tmp[6502]*kernel[1]+tmp[6503]*kernel[2]+tmp[6601]*kernel[3]+tmp[6602]*kernel[4]+tmp[6603]*kernel[5]+tmp[6701]*kernel[6]+tmp[6702]*kernel[7]+tmp[6703]*kernel[8];
				ans[6603]<=tmp[6502]*kernel[0]+tmp[6503]*kernel[1]+tmp[6504]*kernel[2]+tmp[6602]*kernel[3]+tmp[6603]*kernel[4]+tmp[6604]*kernel[5]+tmp[6702]*kernel[6]+tmp[6703]*kernel[7]+tmp[6704]*kernel[8];
				ans[6604]<=tmp[6503]*kernel[0]+tmp[6504]*kernel[1]+tmp[6505]*kernel[2]+tmp[6603]*kernel[3]+tmp[6604]*kernel[4]+tmp[6605]*kernel[5]+tmp[6703]*kernel[6]+tmp[6704]*kernel[7]+tmp[6705]*kernel[8];
				ans[6605]<=tmp[6504]*kernel[0]+tmp[6505]*kernel[1]+tmp[6506]*kernel[2]+tmp[6604]*kernel[3]+tmp[6605]*kernel[4]+tmp[6606]*kernel[5]+tmp[6704]*kernel[6]+tmp[6705]*kernel[7]+tmp[6706]*kernel[8];
				ans[6606]<=tmp[6505]*kernel[0]+tmp[6506]*kernel[1]+tmp[6507]*kernel[2]+tmp[6605]*kernel[3]+tmp[6606]*kernel[4]+tmp[6607]*kernel[5]+tmp[6705]*kernel[6]+tmp[6706]*kernel[7]+tmp[6707]*kernel[8];
				ans[6607]<=tmp[6506]*kernel[0]+tmp[6507]*kernel[1]+tmp[6508]*kernel[2]+tmp[6606]*kernel[3]+tmp[6607]*kernel[4]+tmp[6608]*kernel[5]+tmp[6706]*kernel[6]+tmp[6707]*kernel[7]+tmp[6708]*kernel[8];
				ans[6608]<=tmp[6507]*kernel[0]+tmp[6508]*kernel[1]+tmp[6509]*kernel[2]+tmp[6607]*kernel[3]+tmp[6608]*kernel[4]+tmp[6609]*kernel[5]+tmp[6707]*kernel[6]+tmp[6708]*kernel[7]+tmp[6709]*kernel[8];
				ans[6609]<=tmp[6508]*kernel[0]+tmp[6509]*kernel[1]+tmp[6510]*kernel[2]+tmp[6608]*kernel[3]+tmp[6609]*kernel[4]+tmp[6610]*kernel[5]+tmp[6708]*kernel[6]+tmp[6709]*kernel[7]+tmp[6710]*kernel[8];
				ans[6610]<=tmp[6509]*kernel[0]+tmp[6510]*kernel[1]+tmp[6511]*kernel[2]+tmp[6609]*kernel[3]+tmp[6610]*kernel[4]+tmp[6611]*kernel[5]+tmp[6709]*kernel[6]+tmp[6710]*kernel[7]+tmp[6711]*kernel[8];
				ans[6611]<=tmp[6510]*kernel[0]+tmp[6511]*kernel[1]+tmp[6512]*kernel[2]+tmp[6610]*kernel[3]+tmp[6611]*kernel[4]+tmp[6612]*kernel[5]+tmp[6710]*kernel[6]+tmp[6711]*kernel[7]+tmp[6712]*kernel[8];
				ans[6612]<=tmp[6511]*kernel[0]+tmp[6512]*kernel[1]+tmp[6513]*kernel[2]+tmp[6611]*kernel[3]+tmp[6612]*kernel[4]+tmp[6613]*kernel[5]+tmp[6711]*kernel[6]+tmp[6712]*kernel[7]+tmp[6713]*kernel[8];
				ans[6613]<=tmp[6512]*kernel[0]+tmp[6513]*kernel[1]+tmp[6514]*kernel[2]+tmp[6612]*kernel[3]+tmp[6613]*kernel[4]+tmp[6614]*kernel[5]+tmp[6712]*kernel[6]+tmp[6713]*kernel[7]+tmp[6714]*kernel[8];
				ans[6614]<=tmp[6513]*kernel[0]+tmp[6514]*kernel[1]+tmp[6515]*kernel[2]+tmp[6613]*kernel[3]+tmp[6614]*kernel[4]+tmp[6615]*kernel[5]+tmp[6713]*kernel[6]+tmp[6714]*kernel[7]+tmp[6715]*kernel[8];
				ans[6615]<=tmp[6514]*kernel[0]+tmp[6515]*kernel[1]+tmp[6516]*kernel[2]+tmp[6614]*kernel[3]+tmp[6615]*kernel[4]+tmp[6616]*kernel[5]+tmp[6714]*kernel[6]+tmp[6715]*kernel[7]+tmp[6716]*kernel[8];
				ans[6616]<=tmp[6515]*kernel[0]+tmp[6516]*kernel[1]+tmp[6517]*kernel[2]+tmp[6615]*kernel[3]+tmp[6616]*kernel[4]+tmp[6617]*kernel[5]+tmp[6715]*kernel[6]+tmp[6716]*kernel[7]+tmp[6717]*kernel[8];
				ans[6617]<=tmp[6516]*kernel[0]+tmp[6517]*kernel[1]+tmp[6518]*kernel[2]+tmp[6616]*kernel[3]+tmp[6617]*kernel[4]+tmp[6618]*kernel[5]+tmp[6716]*kernel[6]+tmp[6717]*kernel[7]+tmp[6718]*kernel[8];
				ans[6618]<=tmp[6517]*kernel[0]+tmp[6518]*kernel[1]+tmp[6519]*kernel[2]+tmp[6617]*kernel[3]+tmp[6618]*kernel[4]+tmp[6619]*kernel[5]+tmp[6717]*kernel[6]+tmp[6718]*kernel[7]+tmp[6719]*kernel[8];
				ans[6619]<=tmp[6518]*kernel[0]+tmp[6519]*kernel[1]+tmp[6520]*kernel[2]+tmp[6618]*kernel[3]+tmp[6619]*kernel[4]+tmp[6620]*kernel[5]+tmp[6718]*kernel[6]+tmp[6719]*kernel[7]+tmp[6720]*kernel[8];
				ans[6620]<=tmp[6519]*kernel[0]+tmp[6520]*kernel[1]+tmp[6521]*kernel[2]+tmp[6619]*kernel[3]+tmp[6620]*kernel[4]+tmp[6621]*kernel[5]+tmp[6719]*kernel[6]+tmp[6720]*kernel[7]+tmp[6721]*kernel[8];
				ans[6621]<=tmp[6520]*kernel[0]+tmp[6521]*kernel[1]+tmp[6522]*kernel[2]+tmp[6620]*kernel[3]+tmp[6621]*kernel[4]+tmp[6622]*kernel[5]+tmp[6720]*kernel[6]+tmp[6721]*kernel[7]+tmp[6722]*kernel[8];
				ans[6622]<=tmp[6521]*kernel[0]+tmp[6522]*kernel[1]+tmp[6523]*kernel[2]+tmp[6621]*kernel[3]+tmp[6622]*kernel[4]+tmp[6623]*kernel[5]+tmp[6721]*kernel[6]+tmp[6722]*kernel[7]+tmp[6723]*kernel[8];
				ans[6623]<=tmp[6522]*kernel[0]+tmp[6523]*kernel[1]+tmp[6524]*kernel[2]+tmp[6622]*kernel[3]+tmp[6623]*kernel[4]+tmp[6624]*kernel[5]+tmp[6722]*kernel[6]+tmp[6723]*kernel[7]+tmp[6724]*kernel[8];
				ans[6624]<=tmp[6523]*kernel[0]+tmp[6524]*kernel[1]+tmp[6525]*kernel[2]+tmp[6623]*kernel[3]+tmp[6624]*kernel[4]+tmp[6625]*kernel[5]+tmp[6723]*kernel[6]+tmp[6724]*kernel[7]+tmp[6725]*kernel[8];
				ans[6625]<=tmp[6524]*kernel[0]+tmp[6525]*kernel[1]+tmp[6526]*kernel[2]+tmp[6624]*kernel[3]+tmp[6625]*kernel[4]+tmp[6626]*kernel[5]+tmp[6724]*kernel[6]+tmp[6725]*kernel[7]+tmp[6726]*kernel[8];
				ans[6626]<=tmp[6525]*kernel[0]+tmp[6526]*kernel[1]+tmp[6527]*kernel[2]+tmp[6625]*kernel[3]+tmp[6626]*kernel[4]+tmp[6627]*kernel[5]+tmp[6725]*kernel[6]+tmp[6726]*kernel[7]+tmp[6727]*kernel[8];
				ans[6627]<=tmp[6526]*kernel[0]+tmp[6527]*kernel[1]+tmp[6528]*kernel[2]+tmp[6626]*kernel[3]+tmp[6627]*kernel[4]+tmp[6628]*kernel[5]+tmp[6726]*kernel[6]+tmp[6727]*kernel[7]+tmp[6728]*kernel[8];
				ans[6628]<=tmp[6527]*kernel[0]+tmp[6528]*kernel[1]+tmp[6529]*kernel[2]+tmp[6627]*kernel[3]+tmp[6628]*kernel[4]+tmp[6629]*kernel[5]+tmp[6727]*kernel[6]+tmp[6728]*kernel[7]+tmp[6729]*kernel[8];
				ans[6629]<=tmp[6528]*kernel[0]+tmp[6529]*kernel[1]+tmp[6530]*kernel[2]+tmp[6628]*kernel[3]+tmp[6629]*kernel[4]+tmp[6630]*kernel[5]+tmp[6728]*kernel[6]+tmp[6729]*kernel[7]+tmp[6730]*kernel[8];
				ans[6630]<=tmp[6529]*kernel[0]+tmp[6530]*kernel[1]+tmp[6531]*kernel[2]+tmp[6629]*kernel[3]+tmp[6630]*kernel[4]+tmp[6631]*kernel[5]+tmp[6729]*kernel[6]+tmp[6730]*kernel[7]+tmp[6731]*kernel[8];
				ans[6631]<=tmp[6530]*kernel[0]+tmp[6531]*kernel[1]+tmp[6532]*kernel[2]+tmp[6630]*kernel[3]+tmp[6631]*kernel[4]+tmp[6632]*kernel[5]+tmp[6730]*kernel[6]+tmp[6731]*kernel[7]+tmp[6732]*kernel[8];
				ans[6632]<=tmp[6531]*kernel[0]+tmp[6532]*kernel[1]+tmp[6533]*kernel[2]+tmp[6631]*kernel[3]+tmp[6632]*kernel[4]+tmp[6633]*kernel[5]+tmp[6731]*kernel[6]+tmp[6732]*kernel[7]+tmp[6733]*kernel[8];
				ans[6633]<=tmp[6532]*kernel[0]+tmp[6533]*kernel[1]+tmp[6534]*kernel[2]+tmp[6632]*kernel[3]+tmp[6633]*kernel[4]+tmp[6634]*kernel[5]+tmp[6732]*kernel[6]+tmp[6733]*kernel[7]+tmp[6734]*kernel[8];
				ans[6634]<=tmp[6533]*kernel[0]+tmp[6534]*kernel[1]+tmp[6535]*kernel[2]+tmp[6633]*kernel[3]+tmp[6634]*kernel[4]+tmp[6635]*kernel[5]+tmp[6733]*kernel[6]+tmp[6734]*kernel[7]+tmp[6735]*kernel[8];
				ans[6635]<=tmp[6534]*kernel[0]+tmp[6535]*kernel[1]+tmp[6536]*kernel[2]+tmp[6634]*kernel[3]+tmp[6635]*kernel[4]+tmp[6636]*kernel[5]+tmp[6734]*kernel[6]+tmp[6735]*kernel[7]+tmp[6736]*kernel[8];
				ans[6636]<=tmp[6535]*kernel[0]+tmp[6536]*kernel[1]+tmp[6537]*kernel[2]+tmp[6635]*kernel[3]+tmp[6636]*kernel[4]+tmp[6637]*kernel[5]+tmp[6735]*kernel[6]+tmp[6736]*kernel[7]+tmp[6737]*kernel[8];
				ans[6637]<=tmp[6536]*kernel[0]+tmp[6537]*kernel[1]+tmp[6538]*kernel[2]+tmp[6636]*kernel[3]+tmp[6637]*kernel[4]+tmp[6638]*kernel[5]+tmp[6736]*kernel[6]+tmp[6737]*kernel[7]+tmp[6738]*kernel[8];
				ans[6638]<=tmp[6537]*kernel[0]+tmp[6538]*kernel[1]+tmp[6539]*kernel[2]+tmp[6637]*kernel[3]+tmp[6638]*kernel[4]+tmp[6639]*kernel[5]+tmp[6737]*kernel[6]+tmp[6738]*kernel[7]+tmp[6739]*kernel[8];
				ans[6639]<=tmp[6538]*kernel[0]+tmp[6539]*kernel[1]+tmp[6540]*kernel[2]+tmp[6638]*kernel[3]+tmp[6639]*kernel[4]+tmp[6640]*kernel[5]+tmp[6738]*kernel[6]+tmp[6739]*kernel[7]+tmp[6740]*kernel[8];
				ans[6640]<=tmp[6539]*kernel[0]+tmp[6540]*kernel[1]+tmp[6541]*kernel[2]+tmp[6639]*kernel[3]+tmp[6640]*kernel[4]+tmp[6641]*kernel[5]+tmp[6739]*kernel[6]+tmp[6740]*kernel[7]+tmp[6741]*kernel[8];
				ans[6641]<=tmp[6540]*kernel[0]+tmp[6541]*kernel[1]+tmp[6542]*kernel[2]+tmp[6640]*kernel[3]+tmp[6641]*kernel[4]+tmp[6642]*kernel[5]+tmp[6740]*kernel[6]+tmp[6741]*kernel[7]+tmp[6742]*kernel[8];
				ans[6642]<=tmp[6541]*kernel[0]+tmp[6542]*kernel[1]+tmp[6543]*kernel[2]+tmp[6641]*kernel[3]+tmp[6642]*kernel[4]+tmp[6643]*kernel[5]+tmp[6741]*kernel[6]+tmp[6742]*kernel[7]+tmp[6743]*kernel[8];
				ans[6643]<=tmp[6542]*kernel[0]+tmp[6543]*kernel[1]+tmp[6544]*kernel[2]+tmp[6642]*kernel[3]+tmp[6643]*kernel[4]+tmp[6644]*kernel[5]+tmp[6742]*kernel[6]+tmp[6743]*kernel[7]+tmp[6744]*kernel[8];
				ans[6644]<=tmp[6543]*kernel[0]+tmp[6544]*kernel[1]+tmp[6545]*kernel[2]+tmp[6643]*kernel[3]+tmp[6644]*kernel[4]+tmp[6645]*kernel[5]+tmp[6743]*kernel[6]+tmp[6744]*kernel[7]+tmp[6745]*kernel[8];
				ans[6645]<=tmp[6544]*kernel[0]+tmp[6545]*kernel[1]+tmp[6546]*kernel[2]+tmp[6644]*kernel[3]+tmp[6645]*kernel[4]+tmp[6646]*kernel[5]+tmp[6744]*kernel[6]+tmp[6745]*kernel[7]+tmp[6746]*kernel[8];
				ans[6646]<=tmp[6545]*kernel[0]+tmp[6546]*kernel[1]+tmp[6547]*kernel[2]+tmp[6645]*kernel[3]+tmp[6646]*kernel[4]+tmp[6647]*kernel[5]+tmp[6745]*kernel[6]+tmp[6746]*kernel[7]+tmp[6747]*kernel[8];
				ans[6647]<=tmp[6546]*kernel[0]+tmp[6547]*kernel[1]+tmp[6548]*kernel[2]+tmp[6646]*kernel[3]+tmp[6647]*kernel[4]+tmp[6648]*kernel[5]+tmp[6746]*kernel[6]+tmp[6747]*kernel[7]+tmp[6748]*kernel[8];
				ans[6648]<=tmp[6547]*kernel[0]+tmp[6548]*kernel[1]+tmp[6549]*kernel[2]+tmp[6647]*kernel[3]+tmp[6648]*kernel[4]+tmp[6649]*kernel[5]+tmp[6747]*kernel[6]+tmp[6748]*kernel[7]+tmp[6749]*kernel[8];
				ans[6649]<=tmp[6548]*kernel[0]+tmp[6549]*kernel[1]+tmp[6550]*kernel[2]+tmp[6648]*kernel[3]+tmp[6649]*kernel[4]+tmp[6650]*kernel[5]+tmp[6748]*kernel[6]+tmp[6749]*kernel[7]+tmp[6750]*kernel[8];
				ans[6650]<=tmp[6549]*kernel[0]+tmp[6550]*kernel[1]+tmp[6551]*kernel[2]+tmp[6649]*kernel[3]+tmp[6650]*kernel[4]+tmp[6651]*kernel[5]+tmp[6749]*kernel[6]+tmp[6750]*kernel[7]+tmp[6751]*kernel[8];
				ans[6651]<=tmp[6550]*kernel[0]+tmp[6551]*kernel[1]+tmp[6552]*kernel[2]+tmp[6650]*kernel[3]+tmp[6651]*kernel[4]+tmp[6652]*kernel[5]+tmp[6750]*kernel[6]+tmp[6751]*kernel[7]+tmp[6752]*kernel[8];
				ans[6652]<=tmp[6551]*kernel[0]+tmp[6552]*kernel[1]+tmp[6553]*kernel[2]+tmp[6651]*kernel[3]+tmp[6652]*kernel[4]+tmp[6653]*kernel[5]+tmp[6751]*kernel[6]+tmp[6752]*kernel[7]+tmp[6753]*kernel[8];
				ans[6653]<=tmp[6552]*kernel[0]+tmp[6553]*kernel[1]+tmp[6554]*kernel[2]+tmp[6652]*kernel[3]+tmp[6653]*kernel[4]+tmp[6654]*kernel[5]+tmp[6752]*kernel[6]+tmp[6753]*kernel[7]+tmp[6754]*kernel[8];
				ans[6654]<=tmp[6553]*kernel[0]+tmp[6554]*kernel[1]+tmp[6555]*kernel[2]+tmp[6653]*kernel[3]+tmp[6654]*kernel[4]+tmp[6655]*kernel[5]+tmp[6753]*kernel[6]+tmp[6754]*kernel[7]+tmp[6755]*kernel[8];
				ans[6655]<=tmp[6554]*kernel[0]+tmp[6555]*kernel[1]+tmp[6556]*kernel[2]+tmp[6654]*kernel[3]+tmp[6655]*kernel[4]+tmp[6656]*kernel[5]+tmp[6754]*kernel[6]+tmp[6755]*kernel[7]+tmp[6756]*kernel[8];
				ans[6656]<=tmp[6555]*kernel[0]+tmp[6556]*kernel[1]+tmp[6557]*kernel[2]+tmp[6655]*kernel[3]+tmp[6656]*kernel[4]+tmp[6657]*kernel[5]+tmp[6755]*kernel[6]+tmp[6756]*kernel[7]+tmp[6757]*kernel[8];
				ans[6657]<=tmp[6556]*kernel[0]+tmp[6557]*kernel[1]+tmp[6558]*kernel[2]+tmp[6656]*kernel[3]+tmp[6657]*kernel[4]+tmp[6658]*kernel[5]+tmp[6756]*kernel[6]+tmp[6757]*kernel[7]+tmp[6758]*kernel[8];
				ans[6658]<=tmp[6557]*kernel[0]+tmp[6558]*kernel[1]+tmp[6559]*kernel[2]+tmp[6657]*kernel[3]+tmp[6658]*kernel[4]+tmp[6659]*kernel[5]+tmp[6757]*kernel[6]+tmp[6758]*kernel[7]+tmp[6759]*kernel[8];
				ans[6659]<=tmp[6558]*kernel[0]+tmp[6559]*kernel[1]+tmp[6560]*kernel[2]+tmp[6658]*kernel[3]+tmp[6659]*kernel[4]+tmp[6660]*kernel[5]+tmp[6758]*kernel[6]+tmp[6759]*kernel[7]+tmp[6760]*kernel[8];
				ans[6660]<=tmp[6559]*kernel[0]+tmp[6560]*kernel[1]+tmp[6561]*kernel[2]+tmp[6659]*kernel[3]+tmp[6660]*kernel[4]+tmp[6661]*kernel[5]+tmp[6759]*kernel[6]+tmp[6760]*kernel[7]+tmp[6761]*kernel[8];
				ans[6661]<=tmp[6560]*kernel[0]+tmp[6561]*kernel[1]+tmp[6562]*kernel[2]+tmp[6660]*kernel[3]+tmp[6661]*kernel[4]+tmp[6662]*kernel[5]+tmp[6760]*kernel[6]+tmp[6761]*kernel[7]+tmp[6762]*kernel[8];
				ans[6662]<=tmp[6561]*kernel[0]+tmp[6562]*kernel[1]+tmp[6563]*kernel[2]+tmp[6661]*kernel[3]+tmp[6662]*kernel[4]+tmp[6663]*kernel[5]+tmp[6761]*kernel[6]+tmp[6762]*kernel[7]+tmp[6763]*kernel[8];
				ans[6663]<=tmp[6562]*kernel[0]+tmp[6563]*kernel[1]+tmp[6564]*kernel[2]+tmp[6662]*kernel[3]+tmp[6663]*kernel[4]+tmp[6664]*kernel[5]+tmp[6762]*kernel[6]+tmp[6763]*kernel[7]+tmp[6764]*kernel[8];
				ans[6664]<=tmp[6563]*kernel[0]+tmp[6564]*kernel[1]+tmp[6565]*kernel[2]+tmp[6663]*kernel[3]+tmp[6664]*kernel[4]+tmp[6665]*kernel[5]+tmp[6763]*kernel[6]+tmp[6764]*kernel[7]+tmp[6765]*kernel[8];
				ans[6665]<=tmp[6564]*kernel[0]+tmp[6565]*kernel[1]+tmp[6566]*kernel[2]+tmp[6664]*kernel[3]+tmp[6665]*kernel[4]+tmp[6666]*kernel[5]+tmp[6764]*kernel[6]+tmp[6765]*kernel[7]+tmp[6766]*kernel[8];
				ans[6666]<=tmp[6565]*kernel[0]+tmp[6566]*kernel[1]+tmp[6567]*kernel[2]+tmp[6665]*kernel[3]+tmp[6666]*kernel[4]+tmp[6667]*kernel[5]+tmp[6765]*kernel[6]+tmp[6766]*kernel[7]+tmp[6767]*kernel[8];
				ans[6667]<=tmp[6566]*kernel[0]+tmp[6567]*kernel[1]+tmp[6568]*kernel[2]+tmp[6666]*kernel[3]+tmp[6667]*kernel[4]+tmp[6668]*kernel[5]+tmp[6766]*kernel[6]+tmp[6767]*kernel[7]+tmp[6768]*kernel[8];
				ans[6668]<=tmp[6567]*kernel[0]+tmp[6568]*kernel[1]+tmp[6569]*kernel[2]+tmp[6667]*kernel[3]+tmp[6668]*kernel[4]+tmp[6669]*kernel[5]+tmp[6767]*kernel[6]+tmp[6768]*kernel[7]+tmp[6769]*kernel[8];
				ans[6669]<=tmp[6568]*kernel[0]+tmp[6569]*kernel[1]+tmp[6570]*kernel[2]+tmp[6668]*kernel[3]+tmp[6669]*kernel[4]+tmp[6670]*kernel[5]+tmp[6768]*kernel[6]+tmp[6769]*kernel[7]+tmp[6770]*kernel[8];
				ans[6670]<=tmp[6569]*kernel[0]+tmp[6570]*kernel[1]+tmp[6571]*kernel[2]+tmp[6669]*kernel[3]+tmp[6670]*kernel[4]+tmp[6671]*kernel[5]+tmp[6769]*kernel[6]+tmp[6770]*kernel[7]+tmp[6771]*kernel[8];
				ans[6671]<=tmp[6570]*kernel[0]+tmp[6571]*kernel[1]+tmp[6572]*kernel[2]+tmp[6670]*kernel[3]+tmp[6671]*kernel[4]+tmp[6672]*kernel[5]+tmp[6770]*kernel[6]+tmp[6771]*kernel[7]+tmp[6772]*kernel[8];
				ans[6672]<=tmp[6571]*kernel[0]+tmp[6572]*kernel[1]+tmp[6573]*kernel[2]+tmp[6671]*kernel[3]+tmp[6672]*kernel[4]+tmp[6673]*kernel[5]+tmp[6771]*kernel[6]+tmp[6772]*kernel[7]+tmp[6773]*kernel[8];
				ans[6673]<=tmp[6572]*kernel[0]+tmp[6573]*kernel[1]+tmp[6574]*kernel[2]+tmp[6672]*kernel[3]+tmp[6673]*kernel[4]+tmp[6674]*kernel[5]+tmp[6772]*kernel[6]+tmp[6773]*kernel[7]+tmp[6774]*kernel[8];
				ans[6674]<=tmp[6573]*kernel[0]+tmp[6574]*kernel[1]+tmp[6575]*kernel[2]+tmp[6673]*kernel[3]+tmp[6674]*kernel[4]+tmp[6675]*kernel[5]+tmp[6773]*kernel[6]+tmp[6774]*kernel[7]+tmp[6775]*kernel[8];
				ans[6675]<=tmp[6574]*kernel[0]+tmp[6575]*kernel[1]+tmp[6576]*kernel[2]+tmp[6674]*kernel[3]+tmp[6675]*kernel[4]+tmp[6676]*kernel[5]+tmp[6774]*kernel[6]+tmp[6775]*kernel[7]+tmp[6776]*kernel[8];
				ans[6676]<=tmp[6575]*kernel[0]+tmp[6576]*kernel[1]+tmp[6577]*kernel[2]+tmp[6675]*kernel[3]+tmp[6676]*kernel[4]+tmp[6677]*kernel[5]+tmp[6775]*kernel[6]+tmp[6776]*kernel[7]+tmp[6777]*kernel[8];
				ans[6677]<=tmp[6576]*kernel[0]+tmp[6577]*kernel[1]+tmp[6578]*kernel[2]+tmp[6676]*kernel[3]+tmp[6677]*kernel[4]+tmp[6678]*kernel[5]+tmp[6776]*kernel[6]+tmp[6777]*kernel[7]+tmp[6778]*kernel[8];
				ans[6678]<=tmp[6577]*kernel[0]+tmp[6578]*kernel[1]+tmp[6579]*kernel[2]+tmp[6677]*kernel[3]+tmp[6678]*kernel[4]+tmp[6679]*kernel[5]+tmp[6777]*kernel[6]+tmp[6778]*kernel[7]+tmp[6779]*kernel[8];
				ans[6679]<=tmp[6578]*kernel[0]+tmp[6579]*kernel[1]+tmp[6580]*kernel[2]+tmp[6678]*kernel[3]+tmp[6679]*kernel[4]+tmp[6680]*kernel[5]+tmp[6778]*kernel[6]+tmp[6779]*kernel[7]+tmp[6780]*kernel[8];
				ans[6680]<=tmp[6579]*kernel[0]+tmp[6580]*kernel[1]+tmp[6581]*kernel[2]+tmp[6679]*kernel[3]+tmp[6680]*kernel[4]+tmp[6681]*kernel[5]+tmp[6779]*kernel[6]+tmp[6780]*kernel[7]+tmp[6781]*kernel[8];
				ans[6681]<=tmp[6580]*kernel[0]+tmp[6581]*kernel[1]+tmp[6582]*kernel[2]+tmp[6680]*kernel[3]+tmp[6681]*kernel[4]+tmp[6682]*kernel[5]+tmp[6780]*kernel[6]+tmp[6781]*kernel[7]+tmp[6782]*kernel[8];
				ans[6682]<=tmp[6581]*kernel[0]+tmp[6582]*kernel[1]+tmp[6583]*kernel[2]+tmp[6681]*kernel[3]+tmp[6682]*kernel[4]+tmp[6683]*kernel[5]+tmp[6781]*kernel[6]+tmp[6782]*kernel[7]+tmp[6783]*kernel[8];
				ans[6683]<=tmp[6582]*kernel[0]+tmp[6583]*kernel[1]+tmp[6584]*kernel[2]+tmp[6682]*kernel[3]+tmp[6683]*kernel[4]+tmp[6684]*kernel[5]+tmp[6782]*kernel[6]+tmp[6783]*kernel[7]+tmp[6784]*kernel[8];
				ans[6684]<=tmp[6583]*kernel[0]+tmp[6584]*kernel[1]+tmp[6585]*kernel[2]+tmp[6683]*kernel[3]+tmp[6684]*kernel[4]+tmp[6685]*kernel[5]+tmp[6783]*kernel[6]+tmp[6784]*kernel[7]+tmp[6785]*kernel[8];
				ans[6685]<=tmp[6584]*kernel[0]+tmp[6585]*kernel[1]+tmp[6586]*kernel[2]+tmp[6684]*kernel[3]+tmp[6685]*kernel[4]+tmp[6686]*kernel[5]+tmp[6784]*kernel[6]+tmp[6785]*kernel[7]+tmp[6786]*kernel[8];
				ans[6686]<=tmp[6585]*kernel[0]+tmp[6586]*kernel[1]+tmp[6587]*kernel[2]+tmp[6685]*kernel[3]+tmp[6686]*kernel[4]+tmp[6687]*kernel[5]+tmp[6785]*kernel[6]+tmp[6786]*kernel[7]+tmp[6787]*kernel[8];
				ans[6687]<=tmp[6586]*kernel[0]+tmp[6587]*kernel[1]+tmp[6588]*kernel[2]+tmp[6686]*kernel[3]+tmp[6687]*kernel[4]+tmp[6688]*kernel[5]+tmp[6786]*kernel[6]+tmp[6787]*kernel[7]+tmp[6788]*kernel[8];
				ans[6688]<=tmp[6587]*kernel[0]+tmp[6588]*kernel[1]+tmp[6589]*kernel[2]+tmp[6687]*kernel[3]+tmp[6688]*kernel[4]+tmp[6689]*kernel[5]+tmp[6787]*kernel[6]+tmp[6788]*kernel[7]+tmp[6789]*kernel[8];
				ans[6689]<=tmp[6588]*kernel[0]+tmp[6589]*kernel[1]+tmp[6590]*kernel[2]+tmp[6688]*kernel[3]+tmp[6689]*kernel[4]+tmp[6690]*kernel[5]+tmp[6788]*kernel[6]+tmp[6789]*kernel[7]+tmp[6790]*kernel[8];
				ans[6690]<=tmp[6589]*kernel[0]+tmp[6590]*kernel[1]+tmp[6591]*kernel[2]+tmp[6689]*kernel[3]+tmp[6690]*kernel[4]+tmp[6691]*kernel[5]+tmp[6789]*kernel[6]+tmp[6790]*kernel[7]+tmp[6791]*kernel[8];
				ans[6691]<=tmp[6590]*kernel[0]+tmp[6591]*kernel[1]+tmp[6592]*kernel[2]+tmp[6690]*kernel[3]+tmp[6691]*kernel[4]+tmp[6692]*kernel[5]+tmp[6790]*kernel[6]+tmp[6791]*kernel[7]+tmp[6792]*kernel[8];
				ans[6692]<=tmp[6591]*kernel[0]+tmp[6592]*kernel[1]+tmp[6593]*kernel[2]+tmp[6691]*kernel[3]+tmp[6692]*kernel[4]+tmp[6693]*kernel[5]+tmp[6791]*kernel[6]+tmp[6792]*kernel[7]+tmp[6793]*kernel[8];
				ans[6693]<=tmp[6592]*kernel[0]+tmp[6593]*kernel[1]+tmp[6594]*kernel[2]+tmp[6692]*kernel[3]+tmp[6693]*kernel[4]+tmp[6694]*kernel[5]+tmp[6792]*kernel[6]+tmp[6793]*kernel[7]+tmp[6794]*kernel[8];
				ans[6694]<=tmp[6593]*kernel[0]+tmp[6594]*kernel[1]+tmp[6595]*kernel[2]+tmp[6693]*kernel[3]+tmp[6694]*kernel[4]+tmp[6695]*kernel[5]+tmp[6793]*kernel[6]+tmp[6794]*kernel[7]+tmp[6795]*kernel[8];
				ans[6695]<=tmp[6594]*kernel[0]+tmp[6595]*kernel[1]+tmp[6596]*kernel[2]+tmp[6694]*kernel[3]+tmp[6695]*kernel[4]+tmp[6696]*kernel[5]+tmp[6794]*kernel[6]+tmp[6795]*kernel[7]+tmp[6796]*kernel[8];
				ans[6696]<=tmp[6595]*kernel[0]+tmp[6596]*kernel[1]+tmp[6597]*kernel[2]+tmp[6695]*kernel[3]+tmp[6696]*kernel[4]+tmp[6697]*kernel[5]+tmp[6795]*kernel[6]+tmp[6796]*kernel[7]+tmp[6797]*kernel[8];
				ans[6697]<=tmp[6596]*kernel[0]+tmp[6597]*kernel[1]+tmp[6598]*kernel[2]+tmp[6696]*kernel[3]+tmp[6697]*kernel[4]+tmp[6698]*kernel[5]+tmp[6796]*kernel[6]+tmp[6797]*kernel[7]+tmp[6798]*kernel[8];
				ans[6698]<=tmp[6597]*kernel[0]+tmp[6598]*kernel[1]+tmp[6599]*kernel[2]+tmp[6697]*kernel[3]+tmp[6698]*kernel[4]+tmp[6699]*kernel[5]+tmp[6797]*kernel[6]+tmp[6798]*kernel[7]+tmp[6799]*kernel[8];
				ans[6699]<=tmp[6598]*kernel[0]+tmp[6599]*kernel[1]+tmp[6698]*kernel[3]+tmp[6699]*kernel[4]+tmp[6798]*kernel[6]+tmp[6799]*kernel[7];
				ans[6700]<=tmp[6600]*kernel[1]+tmp[6601]*kernel[2]+tmp[6700]*kernel[4]+tmp[6701]*kernel[5]+tmp[6800]*kernel[7]+tmp[6801]*kernel[8];
				ans[6701]<=tmp[6600]*kernel[0]+tmp[6601]*kernel[1]+tmp[6602]*kernel[2]+tmp[6700]*kernel[3]+tmp[6701]*kernel[4]+tmp[6702]*kernel[5]+tmp[6800]*kernel[6]+tmp[6801]*kernel[7]+tmp[6802]*kernel[8];
				ans[6702]<=tmp[6601]*kernel[0]+tmp[6602]*kernel[1]+tmp[6603]*kernel[2]+tmp[6701]*kernel[3]+tmp[6702]*kernel[4]+tmp[6703]*kernel[5]+tmp[6801]*kernel[6]+tmp[6802]*kernel[7]+tmp[6803]*kernel[8];
				ans[6703]<=tmp[6602]*kernel[0]+tmp[6603]*kernel[1]+tmp[6604]*kernel[2]+tmp[6702]*kernel[3]+tmp[6703]*kernel[4]+tmp[6704]*kernel[5]+tmp[6802]*kernel[6]+tmp[6803]*kernel[7]+tmp[6804]*kernel[8];
				ans[6704]<=tmp[6603]*kernel[0]+tmp[6604]*kernel[1]+tmp[6605]*kernel[2]+tmp[6703]*kernel[3]+tmp[6704]*kernel[4]+tmp[6705]*kernel[5]+tmp[6803]*kernel[6]+tmp[6804]*kernel[7]+tmp[6805]*kernel[8];
				ans[6705]<=tmp[6604]*kernel[0]+tmp[6605]*kernel[1]+tmp[6606]*kernel[2]+tmp[6704]*kernel[3]+tmp[6705]*kernel[4]+tmp[6706]*kernel[5]+tmp[6804]*kernel[6]+tmp[6805]*kernel[7]+tmp[6806]*kernel[8];
				ans[6706]<=tmp[6605]*kernel[0]+tmp[6606]*kernel[1]+tmp[6607]*kernel[2]+tmp[6705]*kernel[3]+tmp[6706]*kernel[4]+tmp[6707]*kernel[5]+tmp[6805]*kernel[6]+tmp[6806]*kernel[7]+tmp[6807]*kernel[8];
				ans[6707]<=tmp[6606]*kernel[0]+tmp[6607]*kernel[1]+tmp[6608]*kernel[2]+tmp[6706]*kernel[3]+tmp[6707]*kernel[4]+tmp[6708]*kernel[5]+tmp[6806]*kernel[6]+tmp[6807]*kernel[7]+tmp[6808]*kernel[8];
				ans[6708]<=tmp[6607]*kernel[0]+tmp[6608]*kernel[1]+tmp[6609]*kernel[2]+tmp[6707]*kernel[3]+tmp[6708]*kernel[4]+tmp[6709]*kernel[5]+tmp[6807]*kernel[6]+tmp[6808]*kernel[7]+tmp[6809]*kernel[8];
				ans[6709]<=tmp[6608]*kernel[0]+tmp[6609]*kernel[1]+tmp[6610]*kernel[2]+tmp[6708]*kernel[3]+tmp[6709]*kernel[4]+tmp[6710]*kernel[5]+tmp[6808]*kernel[6]+tmp[6809]*kernel[7]+tmp[6810]*kernel[8];
				ans[6710]<=tmp[6609]*kernel[0]+tmp[6610]*kernel[1]+tmp[6611]*kernel[2]+tmp[6709]*kernel[3]+tmp[6710]*kernel[4]+tmp[6711]*kernel[5]+tmp[6809]*kernel[6]+tmp[6810]*kernel[7]+tmp[6811]*kernel[8];
				ans[6711]<=tmp[6610]*kernel[0]+tmp[6611]*kernel[1]+tmp[6612]*kernel[2]+tmp[6710]*kernel[3]+tmp[6711]*kernel[4]+tmp[6712]*kernel[5]+tmp[6810]*kernel[6]+tmp[6811]*kernel[7]+tmp[6812]*kernel[8];
				ans[6712]<=tmp[6611]*kernel[0]+tmp[6612]*kernel[1]+tmp[6613]*kernel[2]+tmp[6711]*kernel[3]+tmp[6712]*kernel[4]+tmp[6713]*kernel[5]+tmp[6811]*kernel[6]+tmp[6812]*kernel[7]+tmp[6813]*kernel[8];
				ans[6713]<=tmp[6612]*kernel[0]+tmp[6613]*kernel[1]+tmp[6614]*kernel[2]+tmp[6712]*kernel[3]+tmp[6713]*kernel[4]+tmp[6714]*kernel[5]+tmp[6812]*kernel[6]+tmp[6813]*kernel[7]+tmp[6814]*kernel[8];
				ans[6714]<=tmp[6613]*kernel[0]+tmp[6614]*kernel[1]+tmp[6615]*kernel[2]+tmp[6713]*kernel[3]+tmp[6714]*kernel[4]+tmp[6715]*kernel[5]+tmp[6813]*kernel[6]+tmp[6814]*kernel[7]+tmp[6815]*kernel[8];
				ans[6715]<=tmp[6614]*kernel[0]+tmp[6615]*kernel[1]+tmp[6616]*kernel[2]+tmp[6714]*kernel[3]+tmp[6715]*kernel[4]+tmp[6716]*kernel[5]+tmp[6814]*kernel[6]+tmp[6815]*kernel[7]+tmp[6816]*kernel[8];
				ans[6716]<=tmp[6615]*kernel[0]+tmp[6616]*kernel[1]+tmp[6617]*kernel[2]+tmp[6715]*kernel[3]+tmp[6716]*kernel[4]+tmp[6717]*kernel[5]+tmp[6815]*kernel[6]+tmp[6816]*kernel[7]+tmp[6817]*kernel[8];
				ans[6717]<=tmp[6616]*kernel[0]+tmp[6617]*kernel[1]+tmp[6618]*kernel[2]+tmp[6716]*kernel[3]+tmp[6717]*kernel[4]+tmp[6718]*kernel[5]+tmp[6816]*kernel[6]+tmp[6817]*kernel[7]+tmp[6818]*kernel[8];
				ans[6718]<=tmp[6617]*kernel[0]+tmp[6618]*kernel[1]+tmp[6619]*kernel[2]+tmp[6717]*kernel[3]+tmp[6718]*kernel[4]+tmp[6719]*kernel[5]+tmp[6817]*kernel[6]+tmp[6818]*kernel[7]+tmp[6819]*kernel[8];
				ans[6719]<=tmp[6618]*kernel[0]+tmp[6619]*kernel[1]+tmp[6620]*kernel[2]+tmp[6718]*kernel[3]+tmp[6719]*kernel[4]+tmp[6720]*kernel[5]+tmp[6818]*kernel[6]+tmp[6819]*kernel[7]+tmp[6820]*kernel[8];
				ans[6720]<=tmp[6619]*kernel[0]+tmp[6620]*kernel[1]+tmp[6621]*kernel[2]+tmp[6719]*kernel[3]+tmp[6720]*kernel[4]+tmp[6721]*kernel[5]+tmp[6819]*kernel[6]+tmp[6820]*kernel[7]+tmp[6821]*kernel[8];
				ans[6721]<=tmp[6620]*kernel[0]+tmp[6621]*kernel[1]+tmp[6622]*kernel[2]+tmp[6720]*kernel[3]+tmp[6721]*kernel[4]+tmp[6722]*kernel[5]+tmp[6820]*kernel[6]+tmp[6821]*kernel[7]+tmp[6822]*kernel[8];
				ans[6722]<=tmp[6621]*kernel[0]+tmp[6622]*kernel[1]+tmp[6623]*kernel[2]+tmp[6721]*kernel[3]+tmp[6722]*kernel[4]+tmp[6723]*kernel[5]+tmp[6821]*kernel[6]+tmp[6822]*kernel[7]+tmp[6823]*kernel[8];
				ans[6723]<=tmp[6622]*kernel[0]+tmp[6623]*kernel[1]+tmp[6624]*kernel[2]+tmp[6722]*kernel[3]+tmp[6723]*kernel[4]+tmp[6724]*kernel[5]+tmp[6822]*kernel[6]+tmp[6823]*kernel[7]+tmp[6824]*kernel[8];
				ans[6724]<=tmp[6623]*kernel[0]+tmp[6624]*kernel[1]+tmp[6625]*kernel[2]+tmp[6723]*kernel[3]+tmp[6724]*kernel[4]+tmp[6725]*kernel[5]+tmp[6823]*kernel[6]+tmp[6824]*kernel[7]+tmp[6825]*kernel[8];
				ans[6725]<=tmp[6624]*kernel[0]+tmp[6625]*kernel[1]+tmp[6626]*kernel[2]+tmp[6724]*kernel[3]+tmp[6725]*kernel[4]+tmp[6726]*kernel[5]+tmp[6824]*kernel[6]+tmp[6825]*kernel[7]+tmp[6826]*kernel[8];
				ans[6726]<=tmp[6625]*kernel[0]+tmp[6626]*kernel[1]+tmp[6627]*kernel[2]+tmp[6725]*kernel[3]+tmp[6726]*kernel[4]+tmp[6727]*kernel[5]+tmp[6825]*kernel[6]+tmp[6826]*kernel[7]+tmp[6827]*kernel[8];
				ans[6727]<=tmp[6626]*kernel[0]+tmp[6627]*kernel[1]+tmp[6628]*kernel[2]+tmp[6726]*kernel[3]+tmp[6727]*kernel[4]+tmp[6728]*kernel[5]+tmp[6826]*kernel[6]+tmp[6827]*kernel[7]+tmp[6828]*kernel[8];
				ans[6728]<=tmp[6627]*kernel[0]+tmp[6628]*kernel[1]+tmp[6629]*kernel[2]+tmp[6727]*kernel[3]+tmp[6728]*kernel[4]+tmp[6729]*kernel[5]+tmp[6827]*kernel[6]+tmp[6828]*kernel[7]+tmp[6829]*kernel[8];
				ans[6729]<=tmp[6628]*kernel[0]+tmp[6629]*kernel[1]+tmp[6630]*kernel[2]+tmp[6728]*kernel[3]+tmp[6729]*kernel[4]+tmp[6730]*kernel[5]+tmp[6828]*kernel[6]+tmp[6829]*kernel[7]+tmp[6830]*kernel[8];
				ans[6730]<=tmp[6629]*kernel[0]+tmp[6630]*kernel[1]+tmp[6631]*kernel[2]+tmp[6729]*kernel[3]+tmp[6730]*kernel[4]+tmp[6731]*kernel[5]+tmp[6829]*kernel[6]+tmp[6830]*kernel[7]+tmp[6831]*kernel[8];
				ans[6731]<=tmp[6630]*kernel[0]+tmp[6631]*kernel[1]+tmp[6632]*kernel[2]+tmp[6730]*kernel[3]+tmp[6731]*kernel[4]+tmp[6732]*kernel[5]+tmp[6830]*kernel[6]+tmp[6831]*kernel[7]+tmp[6832]*kernel[8];
				ans[6732]<=tmp[6631]*kernel[0]+tmp[6632]*kernel[1]+tmp[6633]*kernel[2]+tmp[6731]*kernel[3]+tmp[6732]*kernel[4]+tmp[6733]*kernel[5]+tmp[6831]*kernel[6]+tmp[6832]*kernel[7]+tmp[6833]*kernel[8];
				ans[6733]<=tmp[6632]*kernel[0]+tmp[6633]*kernel[1]+tmp[6634]*kernel[2]+tmp[6732]*kernel[3]+tmp[6733]*kernel[4]+tmp[6734]*kernel[5]+tmp[6832]*kernel[6]+tmp[6833]*kernel[7]+tmp[6834]*kernel[8];
				ans[6734]<=tmp[6633]*kernel[0]+tmp[6634]*kernel[1]+tmp[6635]*kernel[2]+tmp[6733]*kernel[3]+tmp[6734]*kernel[4]+tmp[6735]*kernel[5]+tmp[6833]*kernel[6]+tmp[6834]*kernel[7]+tmp[6835]*kernel[8];
				ans[6735]<=tmp[6634]*kernel[0]+tmp[6635]*kernel[1]+tmp[6636]*kernel[2]+tmp[6734]*kernel[3]+tmp[6735]*kernel[4]+tmp[6736]*kernel[5]+tmp[6834]*kernel[6]+tmp[6835]*kernel[7]+tmp[6836]*kernel[8];
				ans[6736]<=tmp[6635]*kernel[0]+tmp[6636]*kernel[1]+tmp[6637]*kernel[2]+tmp[6735]*kernel[3]+tmp[6736]*kernel[4]+tmp[6737]*kernel[5]+tmp[6835]*kernel[6]+tmp[6836]*kernel[7]+tmp[6837]*kernel[8];
				ans[6737]<=tmp[6636]*kernel[0]+tmp[6637]*kernel[1]+tmp[6638]*kernel[2]+tmp[6736]*kernel[3]+tmp[6737]*kernel[4]+tmp[6738]*kernel[5]+tmp[6836]*kernel[6]+tmp[6837]*kernel[7]+tmp[6838]*kernel[8];
				ans[6738]<=tmp[6637]*kernel[0]+tmp[6638]*kernel[1]+tmp[6639]*kernel[2]+tmp[6737]*kernel[3]+tmp[6738]*kernel[4]+tmp[6739]*kernel[5]+tmp[6837]*kernel[6]+tmp[6838]*kernel[7]+tmp[6839]*kernel[8];
				ans[6739]<=tmp[6638]*kernel[0]+tmp[6639]*kernel[1]+tmp[6640]*kernel[2]+tmp[6738]*kernel[3]+tmp[6739]*kernel[4]+tmp[6740]*kernel[5]+tmp[6838]*kernel[6]+tmp[6839]*kernel[7]+tmp[6840]*kernel[8];
				ans[6740]<=tmp[6639]*kernel[0]+tmp[6640]*kernel[1]+tmp[6641]*kernel[2]+tmp[6739]*kernel[3]+tmp[6740]*kernel[4]+tmp[6741]*kernel[5]+tmp[6839]*kernel[6]+tmp[6840]*kernel[7]+tmp[6841]*kernel[8];
				ans[6741]<=tmp[6640]*kernel[0]+tmp[6641]*kernel[1]+tmp[6642]*kernel[2]+tmp[6740]*kernel[3]+tmp[6741]*kernel[4]+tmp[6742]*kernel[5]+tmp[6840]*kernel[6]+tmp[6841]*kernel[7]+tmp[6842]*kernel[8];
				ans[6742]<=tmp[6641]*kernel[0]+tmp[6642]*kernel[1]+tmp[6643]*kernel[2]+tmp[6741]*kernel[3]+tmp[6742]*kernel[4]+tmp[6743]*kernel[5]+tmp[6841]*kernel[6]+tmp[6842]*kernel[7]+tmp[6843]*kernel[8];
				ans[6743]<=tmp[6642]*kernel[0]+tmp[6643]*kernel[1]+tmp[6644]*kernel[2]+tmp[6742]*kernel[3]+tmp[6743]*kernel[4]+tmp[6744]*kernel[5]+tmp[6842]*kernel[6]+tmp[6843]*kernel[7]+tmp[6844]*kernel[8];
				ans[6744]<=tmp[6643]*kernel[0]+tmp[6644]*kernel[1]+tmp[6645]*kernel[2]+tmp[6743]*kernel[3]+tmp[6744]*kernel[4]+tmp[6745]*kernel[5]+tmp[6843]*kernel[6]+tmp[6844]*kernel[7]+tmp[6845]*kernel[8];
				ans[6745]<=tmp[6644]*kernel[0]+tmp[6645]*kernel[1]+tmp[6646]*kernel[2]+tmp[6744]*kernel[3]+tmp[6745]*kernel[4]+tmp[6746]*kernel[5]+tmp[6844]*kernel[6]+tmp[6845]*kernel[7]+tmp[6846]*kernel[8];
				ans[6746]<=tmp[6645]*kernel[0]+tmp[6646]*kernel[1]+tmp[6647]*kernel[2]+tmp[6745]*kernel[3]+tmp[6746]*kernel[4]+tmp[6747]*kernel[5]+tmp[6845]*kernel[6]+tmp[6846]*kernel[7]+tmp[6847]*kernel[8];
				ans[6747]<=tmp[6646]*kernel[0]+tmp[6647]*kernel[1]+tmp[6648]*kernel[2]+tmp[6746]*kernel[3]+tmp[6747]*kernel[4]+tmp[6748]*kernel[5]+tmp[6846]*kernel[6]+tmp[6847]*kernel[7]+tmp[6848]*kernel[8];
				ans[6748]<=tmp[6647]*kernel[0]+tmp[6648]*kernel[1]+tmp[6649]*kernel[2]+tmp[6747]*kernel[3]+tmp[6748]*kernel[4]+tmp[6749]*kernel[5]+tmp[6847]*kernel[6]+tmp[6848]*kernel[7]+tmp[6849]*kernel[8];
				ans[6749]<=tmp[6648]*kernel[0]+tmp[6649]*kernel[1]+tmp[6650]*kernel[2]+tmp[6748]*kernel[3]+tmp[6749]*kernel[4]+tmp[6750]*kernel[5]+tmp[6848]*kernel[6]+tmp[6849]*kernel[7]+tmp[6850]*kernel[8];
				ans[6750]<=tmp[6649]*kernel[0]+tmp[6650]*kernel[1]+tmp[6651]*kernel[2]+tmp[6749]*kernel[3]+tmp[6750]*kernel[4]+tmp[6751]*kernel[5]+tmp[6849]*kernel[6]+tmp[6850]*kernel[7]+tmp[6851]*kernel[8];
				ans[6751]<=tmp[6650]*kernel[0]+tmp[6651]*kernel[1]+tmp[6652]*kernel[2]+tmp[6750]*kernel[3]+tmp[6751]*kernel[4]+tmp[6752]*kernel[5]+tmp[6850]*kernel[6]+tmp[6851]*kernel[7]+tmp[6852]*kernel[8];
				ans[6752]<=tmp[6651]*kernel[0]+tmp[6652]*kernel[1]+tmp[6653]*kernel[2]+tmp[6751]*kernel[3]+tmp[6752]*kernel[4]+tmp[6753]*kernel[5]+tmp[6851]*kernel[6]+tmp[6852]*kernel[7]+tmp[6853]*kernel[8];
				ans[6753]<=tmp[6652]*kernel[0]+tmp[6653]*kernel[1]+tmp[6654]*kernel[2]+tmp[6752]*kernel[3]+tmp[6753]*kernel[4]+tmp[6754]*kernel[5]+tmp[6852]*kernel[6]+tmp[6853]*kernel[7]+tmp[6854]*kernel[8];
				ans[6754]<=tmp[6653]*kernel[0]+tmp[6654]*kernel[1]+tmp[6655]*kernel[2]+tmp[6753]*kernel[3]+tmp[6754]*kernel[4]+tmp[6755]*kernel[5]+tmp[6853]*kernel[6]+tmp[6854]*kernel[7]+tmp[6855]*kernel[8];
				ans[6755]<=tmp[6654]*kernel[0]+tmp[6655]*kernel[1]+tmp[6656]*kernel[2]+tmp[6754]*kernel[3]+tmp[6755]*kernel[4]+tmp[6756]*kernel[5]+tmp[6854]*kernel[6]+tmp[6855]*kernel[7]+tmp[6856]*kernel[8];
				ans[6756]<=tmp[6655]*kernel[0]+tmp[6656]*kernel[1]+tmp[6657]*kernel[2]+tmp[6755]*kernel[3]+tmp[6756]*kernel[4]+tmp[6757]*kernel[5]+tmp[6855]*kernel[6]+tmp[6856]*kernel[7]+tmp[6857]*kernel[8];
				ans[6757]<=tmp[6656]*kernel[0]+tmp[6657]*kernel[1]+tmp[6658]*kernel[2]+tmp[6756]*kernel[3]+tmp[6757]*kernel[4]+tmp[6758]*kernel[5]+tmp[6856]*kernel[6]+tmp[6857]*kernel[7]+tmp[6858]*kernel[8];
				ans[6758]<=tmp[6657]*kernel[0]+tmp[6658]*kernel[1]+tmp[6659]*kernel[2]+tmp[6757]*kernel[3]+tmp[6758]*kernel[4]+tmp[6759]*kernel[5]+tmp[6857]*kernel[6]+tmp[6858]*kernel[7]+tmp[6859]*kernel[8];
				ans[6759]<=tmp[6658]*kernel[0]+tmp[6659]*kernel[1]+tmp[6660]*kernel[2]+tmp[6758]*kernel[3]+tmp[6759]*kernel[4]+tmp[6760]*kernel[5]+tmp[6858]*kernel[6]+tmp[6859]*kernel[7]+tmp[6860]*kernel[8];
				ans[6760]<=tmp[6659]*kernel[0]+tmp[6660]*kernel[1]+tmp[6661]*kernel[2]+tmp[6759]*kernel[3]+tmp[6760]*kernel[4]+tmp[6761]*kernel[5]+tmp[6859]*kernel[6]+tmp[6860]*kernel[7]+tmp[6861]*kernel[8];
				ans[6761]<=tmp[6660]*kernel[0]+tmp[6661]*kernel[1]+tmp[6662]*kernel[2]+tmp[6760]*kernel[3]+tmp[6761]*kernel[4]+tmp[6762]*kernel[5]+tmp[6860]*kernel[6]+tmp[6861]*kernel[7]+tmp[6862]*kernel[8];
				ans[6762]<=tmp[6661]*kernel[0]+tmp[6662]*kernel[1]+tmp[6663]*kernel[2]+tmp[6761]*kernel[3]+tmp[6762]*kernel[4]+tmp[6763]*kernel[5]+tmp[6861]*kernel[6]+tmp[6862]*kernel[7]+tmp[6863]*kernel[8];
				ans[6763]<=tmp[6662]*kernel[0]+tmp[6663]*kernel[1]+tmp[6664]*kernel[2]+tmp[6762]*kernel[3]+tmp[6763]*kernel[4]+tmp[6764]*kernel[5]+tmp[6862]*kernel[6]+tmp[6863]*kernel[7]+tmp[6864]*kernel[8];
				ans[6764]<=tmp[6663]*kernel[0]+tmp[6664]*kernel[1]+tmp[6665]*kernel[2]+tmp[6763]*kernel[3]+tmp[6764]*kernel[4]+tmp[6765]*kernel[5]+tmp[6863]*kernel[6]+tmp[6864]*kernel[7]+tmp[6865]*kernel[8];
				ans[6765]<=tmp[6664]*kernel[0]+tmp[6665]*kernel[1]+tmp[6666]*kernel[2]+tmp[6764]*kernel[3]+tmp[6765]*kernel[4]+tmp[6766]*kernel[5]+tmp[6864]*kernel[6]+tmp[6865]*kernel[7]+tmp[6866]*kernel[8];
				ans[6766]<=tmp[6665]*kernel[0]+tmp[6666]*kernel[1]+tmp[6667]*kernel[2]+tmp[6765]*kernel[3]+tmp[6766]*kernel[4]+tmp[6767]*kernel[5]+tmp[6865]*kernel[6]+tmp[6866]*kernel[7]+tmp[6867]*kernel[8];
				ans[6767]<=tmp[6666]*kernel[0]+tmp[6667]*kernel[1]+tmp[6668]*kernel[2]+tmp[6766]*kernel[3]+tmp[6767]*kernel[4]+tmp[6768]*kernel[5]+tmp[6866]*kernel[6]+tmp[6867]*kernel[7]+tmp[6868]*kernel[8];
				ans[6768]<=tmp[6667]*kernel[0]+tmp[6668]*kernel[1]+tmp[6669]*kernel[2]+tmp[6767]*kernel[3]+tmp[6768]*kernel[4]+tmp[6769]*kernel[5]+tmp[6867]*kernel[6]+tmp[6868]*kernel[7]+tmp[6869]*kernel[8];
				ans[6769]<=tmp[6668]*kernel[0]+tmp[6669]*kernel[1]+tmp[6670]*kernel[2]+tmp[6768]*kernel[3]+tmp[6769]*kernel[4]+tmp[6770]*kernel[5]+tmp[6868]*kernel[6]+tmp[6869]*kernel[7]+tmp[6870]*kernel[8];
				ans[6770]<=tmp[6669]*kernel[0]+tmp[6670]*kernel[1]+tmp[6671]*kernel[2]+tmp[6769]*kernel[3]+tmp[6770]*kernel[4]+tmp[6771]*kernel[5]+tmp[6869]*kernel[6]+tmp[6870]*kernel[7]+tmp[6871]*kernel[8];
				ans[6771]<=tmp[6670]*kernel[0]+tmp[6671]*kernel[1]+tmp[6672]*kernel[2]+tmp[6770]*kernel[3]+tmp[6771]*kernel[4]+tmp[6772]*kernel[5]+tmp[6870]*kernel[6]+tmp[6871]*kernel[7]+tmp[6872]*kernel[8];
				ans[6772]<=tmp[6671]*kernel[0]+tmp[6672]*kernel[1]+tmp[6673]*kernel[2]+tmp[6771]*kernel[3]+tmp[6772]*kernel[4]+tmp[6773]*kernel[5]+tmp[6871]*kernel[6]+tmp[6872]*kernel[7]+tmp[6873]*kernel[8];
				ans[6773]<=tmp[6672]*kernel[0]+tmp[6673]*kernel[1]+tmp[6674]*kernel[2]+tmp[6772]*kernel[3]+tmp[6773]*kernel[4]+tmp[6774]*kernel[5]+tmp[6872]*kernel[6]+tmp[6873]*kernel[7]+tmp[6874]*kernel[8];
				ans[6774]<=tmp[6673]*kernel[0]+tmp[6674]*kernel[1]+tmp[6675]*kernel[2]+tmp[6773]*kernel[3]+tmp[6774]*kernel[4]+tmp[6775]*kernel[5]+tmp[6873]*kernel[6]+tmp[6874]*kernel[7]+tmp[6875]*kernel[8];
				ans[6775]<=tmp[6674]*kernel[0]+tmp[6675]*kernel[1]+tmp[6676]*kernel[2]+tmp[6774]*kernel[3]+tmp[6775]*kernel[4]+tmp[6776]*kernel[5]+tmp[6874]*kernel[6]+tmp[6875]*kernel[7]+tmp[6876]*kernel[8];
				ans[6776]<=tmp[6675]*kernel[0]+tmp[6676]*kernel[1]+tmp[6677]*kernel[2]+tmp[6775]*kernel[3]+tmp[6776]*kernel[4]+tmp[6777]*kernel[5]+tmp[6875]*kernel[6]+tmp[6876]*kernel[7]+tmp[6877]*kernel[8];
				ans[6777]<=tmp[6676]*kernel[0]+tmp[6677]*kernel[1]+tmp[6678]*kernel[2]+tmp[6776]*kernel[3]+tmp[6777]*kernel[4]+tmp[6778]*kernel[5]+tmp[6876]*kernel[6]+tmp[6877]*kernel[7]+tmp[6878]*kernel[8];
				ans[6778]<=tmp[6677]*kernel[0]+tmp[6678]*kernel[1]+tmp[6679]*kernel[2]+tmp[6777]*kernel[3]+tmp[6778]*kernel[4]+tmp[6779]*kernel[5]+tmp[6877]*kernel[6]+tmp[6878]*kernel[7]+tmp[6879]*kernel[8];
				ans[6779]<=tmp[6678]*kernel[0]+tmp[6679]*kernel[1]+tmp[6680]*kernel[2]+tmp[6778]*kernel[3]+tmp[6779]*kernel[4]+tmp[6780]*kernel[5]+tmp[6878]*kernel[6]+tmp[6879]*kernel[7]+tmp[6880]*kernel[8];
				ans[6780]<=tmp[6679]*kernel[0]+tmp[6680]*kernel[1]+tmp[6681]*kernel[2]+tmp[6779]*kernel[3]+tmp[6780]*kernel[4]+tmp[6781]*kernel[5]+tmp[6879]*kernel[6]+tmp[6880]*kernel[7]+tmp[6881]*kernel[8];
				ans[6781]<=tmp[6680]*kernel[0]+tmp[6681]*kernel[1]+tmp[6682]*kernel[2]+tmp[6780]*kernel[3]+tmp[6781]*kernel[4]+tmp[6782]*kernel[5]+tmp[6880]*kernel[6]+tmp[6881]*kernel[7]+tmp[6882]*kernel[8];
				ans[6782]<=tmp[6681]*kernel[0]+tmp[6682]*kernel[1]+tmp[6683]*kernel[2]+tmp[6781]*kernel[3]+tmp[6782]*kernel[4]+tmp[6783]*kernel[5]+tmp[6881]*kernel[6]+tmp[6882]*kernel[7]+tmp[6883]*kernel[8];
				ans[6783]<=tmp[6682]*kernel[0]+tmp[6683]*kernel[1]+tmp[6684]*kernel[2]+tmp[6782]*kernel[3]+tmp[6783]*kernel[4]+tmp[6784]*kernel[5]+tmp[6882]*kernel[6]+tmp[6883]*kernel[7]+tmp[6884]*kernel[8];
				ans[6784]<=tmp[6683]*kernel[0]+tmp[6684]*kernel[1]+tmp[6685]*kernel[2]+tmp[6783]*kernel[3]+tmp[6784]*kernel[4]+tmp[6785]*kernel[5]+tmp[6883]*kernel[6]+tmp[6884]*kernel[7]+tmp[6885]*kernel[8];
				ans[6785]<=tmp[6684]*kernel[0]+tmp[6685]*kernel[1]+tmp[6686]*kernel[2]+tmp[6784]*kernel[3]+tmp[6785]*kernel[4]+tmp[6786]*kernel[5]+tmp[6884]*kernel[6]+tmp[6885]*kernel[7]+tmp[6886]*kernel[8];
				ans[6786]<=tmp[6685]*kernel[0]+tmp[6686]*kernel[1]+tmp[6687]*kernel[2]+tmp[6785]*kernel[3]+tmp[6786]*kernel[4]+tmp[6787]*kernel[5]+tmp[6885]*kernel[6]+tmp[6886]*kernel[7]+tmp[6887]*kernel[8];
				ans[6787]<=tmp[6686]*kernel[0]+tmp[6687]*kernel[1]+tmp[6688]*kernel[2]+tmp[6786]*kernel[3]+tmp[6787]*kernel[4]+tmp[6788]*kernel[5]+tmp[6886]*kernel[6]+tmp[6887]*kernel[7]+tmp[6888]*kernel[8];
				ans[6788]<=tmp[6687]*kernel[0]+tmp[6688]*kernel[1]+tmp[6689]*kernel[2]+tmp[6787]*kernel[3]+tmp[6788]*kernel[4]+tmp[6789]*kernel[5]+tmp[6887]*kernel[6]+tmp[6888]*kernel[7]+tmp[6889]*kernel[8];
				ans[6789]<=tmp[6688]*kernel[0]+tmp[6689]*kernel[1]+tmp[6690]*kernel[2]+tmp[6788]*kernel[3]+tmp[6789]*kernel[4]+tmp[6790]*kernel[5]+tmp[6888]*kernel[6]+tmp[6889]*kernel[7]+tmp[6890]*kernel[8];
				ans[6790]<=tmp[6689]*kernel[0]+tmp[6690]*kernel[1]+tmp[6691]*kernel[2]+tmp[6789]*kernel[3]+tmp[6790]*kernel[4]+tmp[6791]*kernel[5]+tmp[6889]*kernel[6]+tmp[6890]*kernel[7]+tmp[6891]*kernel[8];
				ans[6791]<=tmp[6690]*kernel[0]+tmp[6691]*kernel[1]+tmp[6692]*kernel[2]+tmp[6790]*kernel[3]+tmp[6791]*kernel[4]+tmp[6792]*kernel[5]+tmp[6890]*kernel[6]+tmp[6891]*kernel[7]+tmp[6892]*kernel[8];
				ans[6792]<=tmp[6691]*kernel[0]+tmp[6692]*kernel[1]+tmp[6693]*kernel[2]+tmp[6791]*kernel[3]+tmp[6792]*kernel[4]+tmp[6793]*kernel[5]+tmp[6891]*kernel[6]+tmp[6892]*kernel[7]+tmp[6893]*kernel[8];
				ans[6793]<=tmp[6692]*kernel[0]+tmp[6693]*kernel[1]+tmp[6694]*kernel[2]+tmp[6792]*kernel[3]+tmp[6793]*kernel[4]+tmp[6794]*kernel[5]+tmp[6892]*kernel[6]+tmp[6893]*kernel[7]+tmp[6894]*kernel[8];
				ans[6794]<=tmp[6693]*kernel[0]+tmp[6694]*kernel[1]+tmp[6695]*kernel[2]+tmp[6793]*kernel[3]+tmp[6794]*kernel[4]+tmp[6795]*kernel[5]+tmp[6893]*kernel[6]+tmp[6894]*kernel[7]+tmp[6895]*kernel[8];
				ans[6795]<=tmp[6694]*kernel[0]+tmp[6695]*kernel[1]+tmp[6696]*kernel[2]+tmp[6794]*kernel[3]+tmp[6795]*kernel[4]+tmp[6796]*kernel[5]+tmp[6894]*kernel[6]+tmp[6895]*kernel[7]+tmp[6896]*kernel[8];
				ans[6796]<=tmp[6695]*kernel[0]+tmp[6696]*kernel[1]+tmp[6697]*kernel[2]+tmp[6795]*kernel[3]+tmp[6796]*kernel[4]+tmp[6797]*kernel[5]+tmp[6895]*kernel[6]+tmp[6896]*kernel[7]+tmp[6897]*kernel[8];
				ans[6797]<=tmp[6696]*kernel[0]+tmp[6697]*kernel[1]+tmp[6698]*kernel[2]+tmp[6796]*kernel[3]+tmp[6797]*kernel[4]+tmp[6798]*kernel[5]+tmp[6896]*kernel[6]+tmp[6897]*kernel[7]+tmp[6898]*kernel[8];
				ans[6798]<=tmp[6697]*kernel[0]+tmp[6698]*kernel[1]+tmp[6699]*kernel[2]+tmp[6797]*kernel[3]+tmp[6798]*kernel[4]+tmp[6799]*kernel[5]+tmp[6897]*kernel[6]+tmp[6898]*kernel[7]+tmp[6899]*kernel[8];
				ans[6799]<=tmp[6698]*kernel[0]+tmp[6699]*kernel[1]+tmp[6798]*kernel[3]+tmp[6799]*kernel[4]+tmp[6898]*kernel[6]+tmp[6899]*kernel[7];
				ans[6800]<=tmp[6700]*kernel[1]+tmp[6701]*kernel[2]+tmp[6800]*kernel[4]+tmp[6801]*kernel[5]+tmp[6900]*kernel[7]+tmp[6901]*kernel[8];
				ans[6801]<=tmp[6700]*kernel[0]+tmp[6701]*kernel[1]+tmp[6702]*kernel[2]+tmp[6800]*kernel[3]+tmp[6801]*kernel[4]+tmp[6802]*kernel[5]+tmp[6900]*kernel[6]+tmp[6901]*kernel[7]+tmp[6902]*kernel[8];
				ans[6802]<=tmp[6701]*kernel[0]+tmp[6702]*kernel[1]+tmp[6703]*kernel[2]+tmp[6801]*kernel[3]+tmp[6802]*kernel[4]+tmp[6803]*kernel[5]+tmp[6901]*kernel[6]+tmp[6902]*kernel[7]+tmp[6903]*kernel[8];
				ans[6803]<=tmp[6702]*kernel[0]+tmp[6703]*kernel[1]+tmp[6704]*kernel[2]+tmp[6802]*kernel[3]+tmp[6803]*kernel[4]+tmp[6804]*kernel[5]+tmp[6902]*kernel[6]+tmp[6903]*kernel[7]+tmp[6904]*kernel[8];
				ans[6804]<=tmp[6703]*kernel[0]+tmp[6704]*kernel[1]+tmp[6705]*kernel[2]+tmp[6803]*kernel[3]+tmp[6804]*kernel[4]+tmp[6805]*kernel[5]+tmp[6903]*kernel[6]+tmp[6904]*kernel[7]+tmp[6905]*kernel[8];
				ans[6805]<=tmp[6704]*kernel[0]+tmp[6705]*kernel[1]+tmp[6706]*kernel[2]+tmp[6804]*kernel[3]+tmp[6805]*kernel[4]+tmp[6806]*kernel[5]+tmp[6904]*kernel[6]+tmp[6905]*kernel[7]+tmp[6906]*kernel[8];
				ans[6806]<=tmp[6705]*kernel[0]+tmp[6706]*kernel[1]+tmp[6707]*kernel[2]+tmp[6805]*kernel[3]+tmp[6806]*kernel[4]+tmp[6807]*kernel[5]+tmp[6905]*kernel[6]+tmp[6906]*kernel[7]+tmp[6907]*kernel[8];
				ans[6807]<=tmp[6706]*kernel[0]+tmp[6707]*kernel[1]+tmp[6708]*kernel[2]+tmp[6806]*kernel[3]+tmp[6807]*kernel[4]+tmp[6808]*kernel[5]+tmp[6906]*kernel[6]+tmp[6907]*kernel[7]+tmp[6908]*kernel[8];
				ans[6808]<=tmp[6707]*kernel[0]+tmp[6708]*kernel[1]+tmp[6709]*kernel[2]+tmp[6807]*kernel[3]+tmp[6808]*kernel[4]+tmp[6809]*kernel[5]+tmp[6907]*kernel[6]+tmp[6908]*kernel[7]+tmp[6909]*kernel[8];
				ans[6809]<=tmp[6708]*kernel[0]+tmp[6709]*kernel[1]+tmp[6710]*kernel[2]+tmp[6808]*kernel[3]+tmp[6809]*kernel[4]+tmp[6810]*kernel[5]+tmp[6908]*kernel[6]+tmp[6909]*kernel[7]+tmp[6910]*kernel[8];
				ans[6810]<=tmp[6709]*kernel[0]+tmp[6710]*kernel[1]+tmp[6711]*kernel[2]+tmp[6809]*kernel[3]+tmp[6810]*kernel[4]+tmp[6811]*kernel[5]+tmp[6909]*kernel[6]+tmp[6910]*kernel[7]+tmp[6911]*kernel[8];
				ans[6811]<=tmp[6710]*kernel[0]+tmp[6711]*kernel[1]+tmp[6712]*kernel[2]+tmp[6810]*kernel[3]+tmp[6811]*kernel[4]+tmp[6812]*kernel[5]+tmp[6910]*kernel[6]+tmp[6911]*kernel[7]+tmp[6912]*kernel[8];
				ans[6812]<=tmp[6711]*kernel[0]+tmp[6712]*kernel[1]+tmp[6713]*kernel[2]+tmp[6811]*kernel[3]+tmp[6812]*kernel[4]+tmp[6813]*kernel[5]+tmp[6911]*kernel[6]+tmp[6912]*kernel[7]+tmp[6913]*kernel[8];
				ans[6813]<=tmp[6712]*kernel[0]+tmp[6713]*kernel[1]+tmp[6714]*kernel[2]+tmp[6812]*kernel[3]+tmp[6813]*kernel[4]+tmp[6814]*kernel[5]+tmp[6912]*kernel[6]+tmp[6913]*kernel[7]+tmp[6914]*kernel[8];
				ans[6814]<=tmp[6713]*kernel[0]+tmp[6714]*kernel[1]+tmp[6715]*kernel[2]+tmp[6813]*kernel[3]+tmp[6814]*kernel[4]+tmp[6815]*kernel[5]+tmp[6913]*kernel[6]+tmp[6914]*kernel[7]+tmp[6915]*kernel[8];
				ans[6815]<=tmp[6714]*kernel[0]+tmp[6715]*kernel[1]+tmp[6716]*kernel[2]+tmp[6814]*kernel[3]+tmp[6815]*kernel[4]+tmp[6816]*kernel[5]+tmp[6914]*kernel[6]+tmp[6915]*kernel[7]+tmp[6916]*kernel[8];
				ans[6816]<=tmp[6715]*kernel[0]+tmp[6716]*kernel[1]+tmp[6717]*kernel[2]+tmp[6815]*kernel[3]+tmp[6816]*kernel[4]+tmp[6817]*kernel[5]+tmp[6915]*kernel[6]+tmp[6916]*kernel[7]+tmp[6917]*kernel[8];
				ans[6817]<=tmp[6716]*kernel[0]+tmp[6717]*kernel[1]+tmp[6718]*kernel[2]+tmp[6816]*kernel[3]+tmp[6817]*kernel[4]+tmp[6818]*kernel[5]+tmp[6916]*kernel[6]+tmp[6917]*kernel[7]+tmp[6918]*kernel[8];
				ans[6818]<=tmp[6717]*kernel[0]+tmp[6718]*kernel[1]+tmp[6719]*kernel[2]+tmp[6817]*kernel[3]+tmp[6818]*kernel[4]+tmp[6819]*kernel[5]+tmp[6917]*kernel[6]+tmp[6918]*kernel[7]+tmp[6919]*kernel[8];
				ans[6819]<=tmp[6718]*kernel[0]+tmp[6719]*kernel[1]+tmp[6720]*kernel[2]+tmp[6818]*kernel[3]+tmp[6819]*kernel[4]+tmp[6820]*kernel[5]+tmp[6918]*kernel[6]+tmp[6919]*kernel[7]+tmp[6920]*kernel[8];
				ans[6820]<=tmp[6719]*kernel[0]+tmp[6720]*kernel[1]+tmp[6721]*kernel[2]+tmp[6819]*kernel[3]+tmp[6820]*kernel[4]+tmp[6821]*kernel[5]+tmp[6919]*kernel[6]+tmp[6920]*kernel[7]+tmp[6921]*kernel[8];
				ans[6821]<=tmp[6720]*kernel[0]+tmp[6721]*kernel[1]+tmp[6722]*kernel[2]+tmp[6820]*kernel[3]+tmp[6821]*kernel[4]+tmp[6822]*kernel[5]+tmp[6920]*kernel[6]+tmp[6921]*kernel[7]+tmp[6922]*kernel[8];
				ans[6822]<=tmp[6721]*kernel[0]+tmp[6722]*kernel[1]+tmp[6723]*kernel[2]+tmp[6821]*kernel[3]+tmp[6822]*kernel[4]+tmp[6823]*kernel[5]+tmp[6921]*kernel[6]+tmp[6922]*kernel[7]+tmp[6923]*kernel[8];
				ans[6823]<=tmp[6722]*kernel[0]+tmp[6723]*kernel[1]+tmp[6724]*kernel[2]+tmp[6822]*kernel[3]+tmp[6823]*kernel[4]+tmp[6824]*kernel[5]+tmp[6922]*kernel[6]+tmp[6923]*kernel[7]+tmp[6924]*kernel[8];
				ans[6824]<=tmp[6723]*kernel[0]+tmp[6724]*kernel[1]+tmp[6725]*kernel[2]+tmp[6823]*kernel[3]+tmp[6824]*kernel[4]+tmp[6825]*kernel[5]+tmp[6923]*kernel[6]+tmp[6924]*kernel[7]+tmp[6925]*kernel[8];
				ans[6825]<=tmp[6724]*kernel[0]+tmp[6725]*kernel[1]+tmp[6726]*kernel[2]+tmp[6824]*kernel[3]+tmp[6825]*kernel[4]+tmp[6826]*kernel[5]+tmp[6924]*kernel[6]+tmp[6925]*kernel[7]+tmp[6926]*kernel[8];
				ans[6826]<=tmp[6725]*kernel[0]+tmp[6726]*kernel[1]+tmp[6727]*kernel[2]+tmp[6825]*kernel[3]+tmp[6826]*kernel[4]+tmp[6827]*kernel[5]+tmp[6925]*kernel[6]+tmp[6926]*kernel[7]+tmp[6927]*kernel[8];
				ans[6827]<=tmp[6726]*kernel[0]+tmp[6727]*kernel[1]+tmp[6728]*kernel[2]+tmp[6826]*kernel[3]+tmp[6827]*kernel[4]+tmp[6828]*kernel[5]+tmp[6926]*kernel[6]+tmp[6927]*kernel[7]+tmp[6928]*kernel[8];
				ans[6828]<=tmp[6727]*kernel[0]+tmp[6728]*kernel[1]+tmp[6729]*kernel[2]+tmp[6827]*kernel[3]+tmp[6828]*kernel[4]+tmp[6829]*kernel[5]+tmp[6927]*kernel[6]+tmp[6928]*kernel[7]+tmp[6929]*kernel[8];
				ans[6829]<=tmp[6728]*kernel[0]+tmp[6729]*kernel[1]+tmp[6730]*kernel[2]+tmp[6828]*kernel[3]+tmp[6829]*kernel[4]+tmp[6830]*kernel[5]+tmp[6928]*kernel[6]+tmp[6929]*kernel[7]+tmp[6930]*kernel[8];
				ans[6830]<=tmp[6729]*kernel[0]+tmp[6730]*kernel[1]+tmp[6731]*kernel[2]+tmp[6829]*kernel[3]+tmp[6830]*kernel[4]+tmp[6831]*kernel[5]+tmp[6929]*kernel[6]+tmp[6930]*kernel[7]+tmp[6931]*kernel[8];
				ans[6831]<=tmp[6730]*kernel[0]+tmp[6731]*kernel[1]+tmp[6732]*kernel[2]+tmp[6830]*kernel[3]+tmp[6831]*kernel[4]+tmp[6832]*kernel[5]+tmp[6930]*kernel[6]+tmp[6931]*kernel[7]+tmp[6932]*kernel[8];
				ans[6832]<=tmp[6731]*kernel[0]+tmp[6732]*kernel[1]+tmp[6733]*kernel[2]+tmp[6831]*kernel[3]+tmp[6832]*kernel[4]+tmp[6833]*kernel[5]+tmp[6931]*kernel[6]+tmp[6932]*kernel[7]+tmp[6933]*kernel[8];
				ans[6833]<=tmp[6732]*kernel[0]+tmp[6733]*kernel[1]+tmp[6734]*kernel[2]+tmp[6832]*kernel[3]+tmp[6833]*kernel[4]+tmp[6834]*kernel[5]+tmp[6932]*kernel[6]+tmp[6933]*kernel[7]+tmp[6934]*kernel[8];
				ans[6834]<=tmp[6733]*kernel[0]+tmp[6734]*kernel[1]+tmp[6735]*kernel[2]+tmp[6833]*kernel[3]+tmp[6834]*kernel[4]+tmp[6835]*kernel[5]+tmp[6933]*kernel[6]+tmp[6934]*kernel[7]+tmp[6935]*kernel[8];
				ans[6835]<=tmp[6734]*kernel[0]+tmp[6735]*kernel[1]+tmp[6736]*kernel[2]+tmp[6834]*kernel[3]+tmp[6835]*kernel[4]+tmp[6836]*kernel[5]+tmp[6934]*kernel[6]+tmp[6935]*kernel[7]+tmp[6936]*kernel[8];
				ans[6836]<=tmp[6735]*kernel[0]+tmp[6736]*kernel[1]+tmp[6737]*kernel[2]+tmp[6835]*kernel[3]+tmp[6836]*kernel[4]+tmp[6837]*kernel[5]+tmp[6935]*kernel[6]+tmp[6936]*kernel[7]+tmp[6937]*kernel[8];
				ans[6837]<=tmp[6736]*kernel[0]+tmp[6737]*kernel[1]+tmp[6738]*kernel[2]+tmp[6836]*kernel[3]+tmp[6837]*kernel[4]+tmp[6838]*kernel[5]+tmp[6936]*kernel[6]+tmp[6937]*kernel[7]+tmp[6938]*kernel[8];
				ans[6838]<=tmp[6737]*kernel[0]+tmp[6738]*kernel[1]+tmp[6739]*kernel[2]+tmp[6837]*kernel[3]+tmp[6838]*kernel[4]+tmp[6839]*kernel[5]+tmp[6937]*kernel[6]+tmp[6938]*kernel[7]+tmp[6939]*kernel[8];
				ans[6839]<=tmp[6738]*kernel[0]+tmp[6739]*kernel[1]+tmp[6740]*kernel[2]+tmp[6838]*kernel[3]+tmp[6839]*kernel[4]+tmp[6840]*kernel[5]+tmp[6938]*kernel[6]+tmp[6939]*kernel[7]+tmp[6940]*kernel[8];
				ans[6840]<=tmp[6739]*kernel[0]+tmp[6740]*kernel[1]+tmp[6741]*kernel[2]+tmp[6839]*kernel[3]+tmp[6840]*kernel[4]+tmp[6841]*kernel[5]+tmp[6939]*kernel[6]+tmp[6940]*kernel[7]+tmp[6941]*kernel[8];
				ans[6841]<=tmp[6740]*kernel[0]+tmp[6741]*kernel[1]+tmp[6742]*kernel[2]+tmp[6840]*kernel[3]+tmp[6841]*kernel[4]+tmp[6842]*kernel[5]+tmp[6940]*kernel[6]+tmp[6941]*kernel[7]+tmp[6942]*kernel[8];
				ans[6842]<=tmp[6741]*kernel[0]+tmp[6742]*kernel[1]+tmp[6743]*kernel[2]+tmp[6841]*kernel[3]+tmp[6842]*kernel[4]+tmp[6843]*kernel[5]+tmp[6941]*kernel[6]+tmp[6942]*kernel[7]+tmp[6943]*kernel[8];
				ans[6843]<=tmp[6742]*kernel[0]+tmp[6743]*kernel[1]+tmp[6744]*kernel[2]+tmp[6842]*kernel[3]+tmp[6843]*kernel[4]+tmp[6844]*kernel[5]+tmp[6942]*kernel[6]+tmp[6943]*kernel[7]+tmp[6944]*kernel[8];
				ans[6844]<=tmp[6743]*kernel[0]+tmp[6744]*kernel[1]+tmp[6745]*kernel[2]+tmp[6843]*kernel[3]+tmp[6844]*kernel[4]+tmp[6845]*kernel[5]+tmp[6943]*kernel[6]+tmp[6944]*kernel[7]+tmp[6945]*kernel[8];
				ans[6845]<=tmp[6744]*kernel[0]+tmp[6745]*kernel[1]+tmp[6746]*kernel[2]+tmp[6844]*kernel[3]+tmp[6845]*kernel[4]+tmp[6846]*kernel[5]+tmp[6944]*kernel[6]+tmp[6945]*kernel[7]+tmp[6946]*kernel[8];
				ans[6846]<=tmp[6745]*kernel[0]+tmp[6746]*kernel[1]+tmp[6747]*kernel[2]+tmp[6845]*kernel[3]+tmp[6846]*kernel[4]+tmp[6847]*kernel[5]+tmp[6945]*kernel[6]+tmp[6946]*kernel[7]+tmp[6947]*kernel[8];
				ans[6847]<=tmp[6746]*kernel[0]+tmp[6747]*kernel[1]+tmp[6748]*kernel[2]+tmp[6846]*kernel[3]+tmp[6847]*kernel[4]+tmp[6848]*kernel[5]+tmp[6946]*kernel[6]+tmp[6947]*kernel[7]+tmp[6948]*kernel[8];
				ans[6848]<=tmp[6747]*kernel[0]+tmp[6748]*kernel[1]+tmp[6749]*kernel[2]+tmp[6847]*kernel[3]+tmp[6848]*kernel[4]+tmp[6849]*kernel[5]+tmp[6947]*kernel[6]+tmp[6948]*kernel[7]+tmp[6949]*kernel[8];
				ans[6849]<=tmp[6748]*kernel[0]+tmp[6749]*kernel[1]+tmp[6750]*kernel[2]+tmp[6848]*kernel[3]+tmp[6849]*kernel[4]+tmp[6850]*kernel[5]+tmp[6948]*kernel[6]+tmp[6949]*kernel[7]+tmp[6950]*kernel[8];
				ans[6850]<=tmp[6749]*kernel[0]+tmp[6750]*kernel[1]+tmp[6751]*kernel[2]+tmp[6849]*kernel[3]+tmp[6850]*kernel[4]+tmp[6851]*kernel[5]+tmp[6949]*kernel[6]+tmp[6950]*kernel[7]+tmp[6951]*kernel[8];
				ans[6851]<=tmp[6750]*kernel[0]+tmp[6751]*kernel[1]+tmp[6752]*kernel[2]+tmp[6850]*kernel[3]+tmp[6851]*kernel[4]+tmp[6852]*kernel[5]+tmp[6950]*kernel[6]+tmp[6951]*kernel[7]+tmp[6952]*kernel[8];
				ans[6852]<=tmp[6751]*kernel[0]+tmp[6752]*kernel[1]+tmp[6753]*kernel[2]+tmp[6851]*kernel[3]+tmp[6852]*kernel[4]+tmp[6853]*kernel[5]+tmp[6951]*kernel[6]+tmp[6952]*kernel[7]+tmp[6953]*kernel[8];
				ans[6853]<=tmp[6752]*kernel[0]+tmp[6753]*kernel[1]+tmp[6754]*kernel[2]+tmp[6852]*kernel[3]+tmp[6853]*kernel[4]+tmp[6854]*kernel[5]+tmp[6952]*kernel[6]+tmp[6953]*kernel[7]+tmp[6954]*kernel[8];
				ans[6854]<=tmp[6753]*kernel[0]+tmp[6754]*kernel[1]+tmp[6755]*kernel[2]+tmp[6853]*kernel[3]+tmp[6854]*kernel[4]+tmp[6855]*kernel[5]+tmp[6953]*kernel[6]+tmp[6954]*kernel[7]+tmp[6955]*kernel[8];
				ans[6855]<=tmp[6754]*kernel[0]+tmp[6755]*kernel[1]+tmp[6756]*kernel[2]+tmp[6854]*kernel[3]+tmp[6855]*kernel[4]+tmp[6856]*kernel[5]+tmp[6954]*kernel[6]+tmp[6955]*kernel[7]+tmp[6956]*kernel[8];
				ans[6856]<=tmp[6755]*kernel[0]+tmp[6756]*kernel[1]+tmp[6757]*kernel[2]+tmp[6855]*kernel[3]+tmp[6856]*kernel[4]+tmp[6857]*kernel[5]+tmp[6955]*kernel[6]+tmp[6956]*kernel[7]+tmp[6957]*kernel[8];
				ans[6857]<=tmp[6756]*kernel[0]+tmp[6757]*kernel[1]+tmp[6758]*kernel[2]+tmp[6856]*kernel[3]+tmp[6857]*kernel[4]+tmp[6858]*kernel[5]+tmp[6956]*kernel[6]+tmp[6957]*kernel[7]+tmp[6958]*kernel[8];
				ans[6858]<=tmp[6757]*kernel[0]+tmp[6758]*kernel[1]+tmp[6759]*kernel[2]+tmp[6857]*kernel[3]+tmp[6858]*kernel[4]+tmp[6859]*kernel[5]+tmp[6957]*kernel[6]+tmp[6958]*kernel[7]+tmp[6959]*kernel[8];
				ans[6859]<=tmp[6758]*kernel[0]+tmp[6759]*kernel[1]+tmp[6760]*kernel[2]+tmp[6858]*kernel[3]+tmp[6859]*kernel[4]+tmp[6860]*kernel[5]+tmp[6958]*kernel[6]+tmp[6959]*kernel[7]+tmp[6960]*kernel[8];
				ans[6860]<=tmp[6759]*kernel[0]+tmp[6760]*kernel[1]+tmp[6761]*kernel[2]+tmp[6859]*kernel[3]+tmp[6860]*kernel[4]+tmp[6861]*kernel[5]+tmp[6959]*kernel[6]+tmp[6960]*kernel[7]+tmp[6961]*kernel[8];
				ans[6861]<=tmp[6760]*kernel[0]+tmp[6761]*kernel[1]+tmp[6762]*kernel[2]+tmp[6860]*kernel[3]+tmp[6861]*kernel[4]+tmp[6862]*kernel[5]+tmp[6960]*kernel[6]+tmp[6961]*kernel[7]+tmp[6962]*kernel[8];
				ans[6862]<=tmp[6761]*kernel[0]+tmp[6762]*kernel[1]+tmp[6763]*kernel[2]+tmp[6861]*kernel[3]+tmp[6862]*kernel[4]+tmp[6863]*kernel[5]+tmp[6961]*kernel[6]+tmp[6962]*kernel[7]+tmp[6963]*kernel[8];
				ans[6863]<=tmp[6762]*kernel[0]+tmp[6763]*kernel[1]+tmp[6764]*kernel[2]+tmp[6862]*kernel[3]+tmp[6863]*kernel[4]+tmp[6864]*kernel[5]+tmp[6962]*kernel[6]+tmp[6963]*kernel[7]+tmp[6964]*kernel[8];
				ans[6864]<=tmp[6763]*kernel[0]+tmp[6764]*kernel[1]+tmp[6765]*kernel[2]+tmp[6863]*kernel[3]+tmp[6864]*kernel[4]+tmp[6865]*kernel[5]+tmp[6963]*kernel[6]+tmp[6964]*kernel[7]+tmp[6965]*kernel[8];
				ans[6865]<=tmp[6764]*kernel[0]+tmp[6765]*kernel[1]+tmp[6766]*kernel[2]+tmp[6864]*kernel[3]+tmp[6865]*kernel[4]+tmp[6866]*kernel[5]+tmp[6964]*kernel[6]+tmp[6965]*kernel[7]+tmp[6966]*kernel[8];
				ans[6866]<=tmp[6765]*kernel[0]+tmp[6766]*kernel[1]+tmp[6767]*kernel[2]+tmp[6865]*kernel[3]+tmp[6866]*kernel[4]+tmp[6867]*kernel[5]+tmp[6965]*kernel[6]+tmp[6966]*kernel[7]+tmp[6967]*kernel[8];
				ans[6867]<=tmp[6766]*kernel[0]+tmp[6767]*kernel[1]+tmp[6768]*kernel[2]+tmp[6866]*kernel[3]+tmp[6867]*kernel[4]+tmp[6868]*kernel[5]+tmp[6966]*kernel[6]+tmp[6967]*kernel[7]+tmp[6968]*kernel[8];
				ans[6868]<=tmp[6767]*kernel[0]+tmp[6768]*kernel[1]+tmp[6769]*kernel[2]+tmp[6867]*kernel[3]+tmp[6868]*kernel[4]+tmp[6869]*kernel[5]+tmp[6967]*kernel[6]+tmp[6968]*kernel[7]+tmp[6969]*kernel[8];
				ans[6869]<=tmp[6768]*kernel[0]+tmp[6769]*kernel[1]+tmp[6770]*kernel[2]+tmp[6868]*kernel[3]+tmp[6869]*kernel[4]+tmp[6870]*kernel[5]+tmp[6968]*kernel[6]+tmp[6969]*kernel[7]+tmp[6970]*kernel[8];
				ans[6870]<=tmp[6769]*kernel[0]+tmp[6770]*kernel[1]+tmp[6771]*kernel[2]+tmp[6869]*kernel[3]+tmp[6870]*kernel[4]+tmp[6871]*kernel[5]+tmp[6969]*kernel[6]+tmp[6970]*kernel[7]+tmp[6971]*kernel[8];
				ans[6871]<=tmp[6770]*kernel[0]+tmp[6771]*kernel[1]+tmp[6772]*kernel[2]+tmp[6870]*kernel[3]+tmp[6871]*kernel[4]+tmp[6872]*kernel[5]+tmp[6970]*kernel[6]+tmp[6971]*kernel[7]+tmp[6972]*kernel[8];
				ans[6872]<=tmp[6771]*kernel[0]+tmp[6772]*kernel[1]+tmp[6773]*kernel[2]+tmp[6871]*kernel[3]+tmp[6872]*kernel[4]+tmp[6873]*kernel[5]+tmp[6971]*kernel[6]+tmp[6972]*kernel[7]+tmp[6973]*kernel[8];
				ans[6873]<=tmp[6772]*kernel[0]+tmp[6773]*kernel[1]+tmp[6774]*kernel[2]+tmp[6872]*kernel[3]+tmp[6873]*kernel[4]+tmp[6874]*kernel[5]+tmp[6972]*kernel[6]+tmp[6973]*kernel[7]+tmp[6974]*kernel[8];
				ans[6874]<=tmp[6773]*kernel[0]+tmp[6774]*kernel[1]+tmp[6775]*kernel[2]+tmp[6873]*kernel[3]+tmp[6874]*kernel[4]+tmp[6875]*kernel[5]+tmp[6973]*kernel[6]+tmp[6974]*kernel[7]+tmp[6975]*kernel[8];
				ans[6875]<=tmp[6774]*kernel[0]+tmp[6775]*kernel[1]+tmp[6776]*kernel[2]+tmp[6874]*kernel[3]+tmp[6875]*kernel[4]+tmp[6876]*kernel[5]+tmp[6974]*kernel[6]+tmp[6975]*kernel[7]+tmp[6976]*kernel[8];
				ans[6876]<=tmp[6775]*kernel[0]+tmp[6776]*kernel[1]+tmp[6777]*kernel[2]+tmp[6875]*kernel[3]+tmp[6876]*kernel[4]+tmp[6877]*kernel[5]+tmp[6975]*kernel[6]+tmp[6976]*kernel[7]+tmp[6977]*kernel[8];
				ans[6877]<=tmp[6776]*kernel[0]+tmp[6777]*kernel[1]+tmp[6778]*kernel[2]+tmp[6876]*kernel[3]+tmp[6877]*kernel[4]+tmp[6878]*kernel[5]+tmp[6976]*kernel[6]+tmp[6977]*kernel[7]+tmp[6978]*kernel[8];
				ans[6878]<=tmp[6777]*kernel[0]+tmp[6778]*kernel[1]+tmp[6779]*kernel[2]+tmp[6877]*kernel[3]+tmp[6878]*kernel[4]+tmp[6879]*kernel[5]+tmp[6977]*kernel[6]+tmp[6978]*kernel[7]+tmp[6979]*kernel[8];
				ans[6879]<=tmp[6778]*kernel[0]+tmp[6779]*kernel[1]+tmp[6780]*kernel[2]+tmp[6878]*kernel[3]+tmp[6879]*kernel[4]+tmp[6880]*kernel[5]+tmp[6978]*kernel[6]+tmp[6979]*kernel[7]+tmp[6980]*kernel[8];
				ans[6880]<=tmp[6779]*kernel[0]+tmp[6780]*kernel[1]+tmp[6781]*kernel[2]+tmp[6879]*kernel[3]+tmp[6880]*kernel[4]+tmp[6881]*kernel[5]+tmp[6979]*kernel[6]+tmp[6980]*kernel[7]+tmp[6981]*kernel[8];
				ans[6881]<=tmp[6780]*kernel[0]+tmp[6781]*kernel[1]+tmp[6782]*kernel[2]+tmp[6880]*kernel[3]+tmp[6881]*kernel[4]+tmp[6882]*kernel[5]+tmp[6980]*kernel[6]+tmp[6981]*kernel[7]+tmp[6982]*kernel[8];
				ans[6882]<=tmp[6781]*kernel[0]+tmp[6782]*kernel[1]+tmp[6783]*kernel[2]+tmp[6881]*kernel[3]+tmp[6882]*kernel[4]+tmp[6883]*kernel[5]+tmp[6981]*kernel[6]+tmp[6982]*kernel[7]+tmp[6983]*kernel[8];
				ans[6883]<=tmp[6782]*kernel[0]+tmp[6783]*kernel[1]+tmp[6784]*kernel[2]+tmp[6882]*kernel[3]+tmp[6883]*kernel[4]+tmp[6884]*kernel[5]+tmp[6982]*kernel[6]+tmp[6983]*kernel[7]+tmp[6984]*kernel[8];
				ans[6884]<=tmp[6783]*kernel[0]+tmp[6784]*kernel[1]+tmp[6785]*kernel[2]+tmp[6883]*kernel[3]+tmp[6884]*kernel[4]+tmp[6885]*kernel[5]+tmp[6983]*kernel[6]+tmp[6984]*kernel[7]+tmp[6985]*kernel[8];
				ans[6885]<=tmp[6784]*kernel[0]+tmp[6785]*kernel[1]+tmp[6786]*kernel[2]+tmp[6884]*kernel[3]+tmp[6885]*kernel[4]+tmp[6886]*kernel[5]+tmp[6984]*kernel[6]+tmp[6985]*kernel[7]+tmp[6986]*kernel[8];
				ans[6886]<=tmp[6785]*kernel[0]+tmp[6786]*kernel[1]+tmp[6787]*kernel[2]+tmp[6885]*kernel[3]+tmp[6886]*kernel[4]+tmp[6887]*kernel[5]+tmp[6985]*kernel[6]+tmp[6986]*kernel[7]+tmp[6987]*kernel[8];
				ans[6887]<=tmp[6786]*kernel[0]+tmp[6787]*kernel[1]+tmp[6788]*kernel[2]+tmp[6886]*kernel[3]+tmp[6887]*kernel[4]+tmp[6888]*kernel[5]+tmp[6986]*kernel[6]+tmp[6987]*kernel[7]+tmp[6988]*kernel[8];
				ans[6888]<=tmp[6787]*kernel[0]+tmp[6788]*kernel[1]+tmp[6789]*kernel[2]+tmp[6887]*kernel[3]+tmp[6888]*kernel[4]+tmp[6889]*kernel[5]+tmp[6987]*kernel[6]+tmp[6988]*kernel[7]+tmp[6989]*kernel[8];
				ans[6889]<=tmp[6788]*kernel[0]+tmp[6789]*kernel[1]+tmp[6790]*kernel[2]+tmp[6888]*kernel[3]+tmp[6889]*kernel[4]+tmp[6890]*kernel[5]+tmp[6988]*kernel[6]+tmp[6989]*kernel[7]+tmp[6990]*kernel[8];
				ans[6890]<=tmp[6789]*kernel[0]+tmp[6790]*kernel[1]+tmp[6791]*kernel[2]+tmp[6889]*kernel[3]+tmp[6890]*kernel[4]+tmp[6891]*kernel[5]+tmp[6989]*kernel[6]+tmp[6990]*kernel[7]+tmp[6991]*kernel[8];
				ans[6891]<=tmp[6790]*kernel[0]+tmp[6791]*kernel[1]+tmp[6792]*kernel[2]+tmp[6890]*kernel[3]+tmp[6891]*kernel[4]+tmp[6892]*kernel[5]+tmp[6990]*kernel[6]+tmp[6991]*kernel[7]+tmp[6992]*kernel[8];
				ans[6892]<=tmp[6791]*kernel[0]+tmp[6792]*kernel[1]+tmp[6793]*kernel[2]+tmp[6891]*kernel[3]+tmp[6892]*kernel[4]+tmp[6893]*kernel[5]+tmp[6991]*kernel[6]+tmp[6992]*kernel[7]+tmp[6993]*kernel[8];
				ans[6893]<=tmp[6792]*kernel[0]+tmp[6793]*kernel[1]+tmp[6794]*kernel[2]+tmp[6892]*kernel[3]+tmp[6893]*kernel[4]+tmp[6894]*kernel[5]+tmp[6992]*kernel[6]+tmp[6993]*kernel[7]+tmp[6994]*kernel[8];
				ans[6894]<=tmp[6793]*kernel[0]+tmp[6794]*kernel[1]+tmp[6795]*kernel[2]+tmp[6893]*kernel[3]+tmp[6894]*kernel[4]+tmp[6895]*kernel[5]+tmp[6993]*kernel[6]+tmp[6994]*kernel[7]+tmp[6995]*kernel[8];
				ans[6895]<=tmp[6794]*kernel[0]+tmp[6795]*kernel[1]+tmp[6796]*kernel[2]+tmp[6894]*kernel[3]+tmp[6895]*kernel[4]+tmp[6896]*kernel[5]+tmp[6994]*kernel[6]+tmp[6995]*kernel[7]+tmp[6996]*kernel[8];
				ans[6896]<=tmp[6795]*kernel[0]+tmp[6796]*kernel[1]+tmp[6797]*kernel[2]+tmp[6895]*kernel[3]+tmp[6896]*kernel[4]+tmp[6897]*kernel[5]+tmp[6995]*kernel[6]+tmp[6996]*kernel[7]+tmp[6997]*kernel[8];
				ans[6897]<=tmp[6796]*kernel[0]+tmp[6797]*kernel[1]+tmp[6798]*kernel[2]+tmp[6896]*kernel[3]+tmp[6897]*kernel[4]+tmp[6898]*kernel[5]+tmp[6996]*kernel[6]+tmp[6997]*kernel[7]+tmp[6998]*kernel[8];
				ans[6898]<=tmp[6797]*kernel[0]+tmp[6798]*kernel[1]+tmp[6799]*kernel[2]+tmp[6897]*kernel[3]+tmp[6898]*kernel[4]+tmp[6899]*kernel[5]+tmp[6997]*kernel[6]+tmp[6998]*kernel[7]+tmp[6999]*kernel[8];
				ans[6899]<=tmp[6798]*kernel[0]+tmp[6799]*kernel[1]+tmp[6898]*kernel[3]+tmp[6899]*kernel[4]+tmp[6998]*kernel[6]+tmp[6999]*kernel[7];
				ans[6900]<=tmp[6800]*kernel[1]+tmp[6801]*kernel[2]+tmp[6900]*kernel[4]+tmp[6901]*kernel[5]+tmp[7000]*kernel[7]+tmp[7001]*kernel[8];
				ans[6901]<=tmp[6800]*kernel[0]+tmp[6801]*kernel[1]+tmp[6802]*kernel[2]+tmp[6900]*kernel[3]+tmp[6901]*kernel[4]+tmp[6902]*kernel[5]+tmp[7000]*kernel[6]+tmp[7001]*kernel[7]+tmp[7002]*kernel[8];
				ans[6902]<=tmp[6801]*kernel[0]+tmp[6802]*kernel[1]+tmp[6803]*kernel[2]+tmp[6901]*kernel[3]+tmp[6902]*kernel[4]+tmp[6903]*kernel[5]+tmp[7001]*kernel[6]+tmp[7002]*kernel[7]+tmp[7003]*kernel[8];
				ans[6903]<=tmp[6802]*kernel[0]+tmp[6803]*kernel[1]+tmp[6804]*kernel[2]+tmp[6902]*kernel[3]+tmp[6903]*kernel[4]+tmp[6904]*kernel[5]+tmp[7002]*kernel[6]+tmp[7003]*kernel[7]+tmp[7004]*kernel[8];
				ans[6904]<=tmp[6803]*kernel[0]+tmp[6804]*kernel[1]+tmp[6805]*kernel[2]+tmp[6903]*kernel[3]+tmp[6904]*kernel[4]+tmp[6905]*kernel[5]+tmp[7003]*kernel[6]+tmp[7004]*kernel[7]+tmp[7005]*kernel[8];
				ans[6905]<=tmp[6804]*kernel[0]+tmp[6805]*kernel[1]+tmp[6806]*kernel[2]+tmp[6904]*kernel[3]+tmp[6905]*kernel[4]+tmp[6906]*kernel[5]+tmp[7004]*kernel[6]+tmp[7005]*kernel[7]+tmp[7006]*kernel[8];
				ans[6906]<=tmp[6805]*kernel[0]+tmp[6806]*kernel[1]+tmp[6807]*kernel[2]+tmp[6905]*kernel[3]+tmp[6906]*kernel[4]+tmp[6907]*kernel[5]+tmp[7005]*kernel[6]+tmp[7006]*kernel[7]+tmp[7007]*kernel[8];
				ans[6907]<=tmp[6806]*kernel[0]+tmp[6807]*kernel[1]+tmp[6808]*kernel[2]+tmp[6906]*kernel[3]+tmp[6907]*kernel[4]+tmp[6908]*kernel[5]+tmp[7006]*kernel[6]+tmp[7007]*kernel[7]+tmp[7008]*kernel[8];
				ans[6908]<=tmp[6807]*kernel[0]+tmp[6808]*kernel[1]+tmp[6809]*kernel[2]+tmp[6907]*kernel[3]+tmp[6908]*kernel[4]+tmp[6909]*kernel[5]+tmp[7007]*kernel[6]+tmp[7008]*kernel[7]+tmp[7009]*kernel[8];
				ans[6909]<=tmp[6808]*kernel[0]+tmp[6809]*kernel[1]+tmp[6810]*kernel[2]+tmp[6908]*kernel[3]+tmp[6909]*kernel[4]+tmp[6910]*kernel[5]+tmp[7008]*kernel[6]+tmp[7009]*kernel[7]+tmp[7010]*kernel[8];
				ans[6910]<=tmp[6809]*kernel[0]+tmp[6810]*kernel[1]+tmp[6811]*kernel[2]+tmp[6909]*kernel[3]+tmp[6910]*kernel[4]+tmp[6911]*kernel[5]+tmp[7009]*kernel[6]+tmp[7010]*kernel[7]+tmp[7011]*kernel[8];
				ans[6911]<=tmp[6810]*kernel[0]+tmp[6811]*kernel[1]+tmp[6812]*kernel[2]+tmp[6910]*kernel[3]+tmp[6911]*kernel[4]+tmp[6912]*kernel[5]+tmp[7010]*kernel[6]+tmp[7011]*kernel[7]+tmp[7012]*kernel[8];
				ans[6912]<=tmp[6811]*kernel[0]+tmp[6812]*kernel[1]+tmp[6813]*kernel[2]+tmp[6911]*kernel[3]+tmp[6912]*kernel[4]+tmp[6913]*kernel[5]+tmp[7011]*kernel[6]+tmp[7012]*kernel[7]+tmp[7013]*kernel[8];
				ans[6913]<=tmp[6812]*kernel[0]+tmp[6813]*kernel[1]+tmp[6814]*kernel[2]+tmp[6912]*kernel[3]+tmp[6913]*kernel[4]+tmp[6914]*kernel[5]+tmp[7012]*kernel[6]+tmp[7013]*kernel[7]+tmp[7014]*kernel[8];
				ans[6914]<=tmp[6813]*kernel[0]+tmp[6814]*kernel[1]+tmp[6815]*kernel[2]+tmp[6913]*kernel[3]+tmp[6914]*kernel[4]+tmp[6915]*kernel[5]+tmp[7013]*kernel[6]+tmp[7014]*kernel[7]+tmp[7015]*kernel[8];
				ans[6915]<=tmp[6814]*kernel[0]+tmp[6815]*kernel[1]+tmp[6816]*kernel[2]+tmp[6914]*kernel[3]+tmp[6915]*kernel[4]+tmp[6916]*kernel[5]+tmp[7014]*kernel[6]+tmp[7015]*kernel[7]+tmp[7016]*kernel[8];
				ans[6916]<=tmp[6815]*kernel[0]+tmp[6816]*kernel[1]+tmp[6817]*kernel[2]+tmp[6915]*kernel[3]+tmp[6916]*kernel[4]+tmp[6917]*kernel[5]+tmp[7015]*kernel[6]+tmp[7016]*kernel[7]+tmp[7017]*kernel[8];
				ans[6917]<=tmp[6816]*kernel[0]+tmp[6817]*kernel[1]+tmp[6818]*kernel[2]+tmp[6916]*kernel[3]+tmp[6917]*kernel[4]+tmp[6918]*kernel[5]+tmp[7016]*kernel[6]+tmp[7017]*kernel[7]+tmp[7018]*kernel[8];
				ans[6918]<=tmp[6817]*kernel[0]+tmp[6818]*kernel[1]+tmp[6819]*kernel[2]+tmp[6917]*kernel[3]+tmp[6918]*kernel[4]+tmp[6919]*kernel[5]+tmp[7017]*kernel[6]+tmp[7018]*kernel[7]+tmp[7019]*kernel[8];
				ans[6919]<=tmp[6818]*kernel[0]+tmp[6819]*kernel[1]+tmp[6820]*kernel[2]+tmp[6918]*kernel[3]+tmp[6919]*kernel[4]+tmp[6920]*kernel[5]+tmp[7018]*kernel[6]+tmp[7019]*kernel[7]+tmp[7020]*kernel[8];
				ans[6920]<=tmp[6819]*kernel[0]+tmp[6820]*kernel[1]+tmp[6821]*kernel[2]+tmp[6919]*kernel[3]+tmp[6920]*kernel[4]+tmp[6921]*kernel[5]+tmp[7019]*kernel[6]+tmp[7020]*kernel[7]+tmp[7021]*kernel[8];
				ans[6921]<=tmp[6820]*kernel[0]+tmp[6821]*kernel[1]+tmp[6822]*kernel[2]+tmp[6920]*kernel[3]+tmp[6921]*kernel[4]+tmp[6922]*kernel[5]+tmp[7020]*kernel[6]+tmp[7021]*kernel[7]+tmp[7022]*kernel[8];
				ans[6922]<=tmp[6821]*kernel[0]+tmp[6822]*kernel[1]+tmp[6823]*kernel[2]+tmp[6921]*kernel[3]+tmp[6922]*kernel[4]+tmp[6923]*kernel[5]+tmp[7021]*kernel[6]+tmp[7022]*kernel[7]+tmp[7023]*kernel[8];
				ans[6923]<=tmp[6822]*kernel[0]+tmp[6823]*kernel[1]+tmp[6824]*kernel[2]+tmp[6922]*kernel[3]+tmp[6923]*kernel[4]+tmp[6924]*kernel[5]+tmp[7022]*kernel[6]+tmp[7023]*kernel[7]+tmp[7024]*kernel[8];
				ans[6924]<=tmp[6823]*kernel[0]+tmp[6824]*kernel[1]+tmp[6825]*kernel[2]+tmp[6923]*kernel[3]+tmp[6924]*kernel[4]+tmp[6925]*kernel[5]+tmp[7023]*kernel[6]+tmp[7024]*kernel[7]+tmp[7025]*kernel[8];
				ans[6925]<=tmp[6824]*kernel[0]+tmp[6825]*kernel[1]+tmp[6826]*kernel[2]+tmp[6924]*kernel[3]+tmp[6925]*kernel[4]+tmp[6926]*kernel[5]+tmp[7024]*kernel[6]+tmp[7025]*kernel[7]+tmp[7026]*kernel[8];
				ans[6926]<=tmp[6825]*kernel[0]+tmp[6826]*kernel[1]+tmp[6827]*kernel[2]+tmp[6925]*kernel[3]+tmp[6926]*kernel[4]+tmp[6927]*kernel[5]+tmp[7025]*kernel[6]+tmp[7026]*kernel[7]+tmp[7027]*kernel[8];
				ans[6927]<=tmp[6826]*kernel[0]+tmp[6827]*kernel[1]+tmp[6828]*kernel[2]+tmp[6926]*kernel[3]+tmp[6927]*kernel[4]+tmp[6928]*kernel[5]+tmp[7026]*kernel[6]+tmp[7027]*kernel[7]+tmp[7028]*kernel[8];
				ans[6928]<=tmp[6827]*kernel[0]+tmp[6828]*kernel[1]+tmp[6829]*kernel[2]+tmp[6927]*kernel[3]+tmp[6928]*kernel[4]+tmp[6929]*kernel[5]+tmp[7027]*kernel[6]+tmp[7028]*kernel[7]+tmp[7029]*kernel[8];
				ans[6929]<=tmp[6828]*kernel[0]+tmp[6829]*kernel[1]+tmp[6830]*kernel[2]+tmp[6928]*kernel[3]+tmp[6929]*kernel[4]+tmp[6930]*kernel[5]+tmp[7028]*kernel[6]+tmp[7029]*kernel[7]+tmp[7030]*kernel[8];
				ans[6930]<=tmp[6829]*kernel[0]+tmp[6830]*kernel[1]+tmp[6831]*kernel[2]+tmp[6929]*kernel[3]+tmp[6930]*kernel[4]+tmp[6931]*kernel[5]+tmp[7029]*kernel[6]+tmp[7030]*kernel[7]+tmp[7031]*kernel[8];
				ans[6931]<=tmp[6830]*kernel[0]+tmp[6831]*kernel[1]+tmp[6832]*kernel[2]+tmp[6930]*kernel[3]+tmp[6931]*kernel[4]+tmp[6932]*kernel[5]+tmp[7030]*kernel[6]+tmp[7031]*kernel[7]+tmp[7032]*kernel[8];
				ans[6932]<=tmp[6831]*kernel[0]+tmp[6832]*kernel[1]+tmp[6833]*kernel[2]+tmp[6931]*kernel[3]+tmp[6932]*kernel[4]+tmp[6933]*kernel[5]+tmp[7031]*kernel[6]+tmp[7032]*kernel[7]+tmp[7033]*kernel[8];
				ans[6933]<=tmp[6832]*kernel[0]+tmp[6833]*kernel[1]+tmp[6834]*kernel[2]+tmp[6932]*kernel[3]+tmp[6933]*kernel[4]+tmp[6934]*kernel[5]+tmp[7032]*kernel[6]+tmp[7033]*kernel[7]+tmp[7034]*kernel[8];
				ans[6934]<=tmp[6833]*kernel[0]+tmp[6834]*kernel[1]+tmp[6835]*kernel[2]+tmp[6933]*kernel[3]+tmp[6934]*kernel[4]+tmp[6935]*kernel[5]+tmp[7033]*kernel[6]+tmp[7034]*kernel[7]+tmp[7035]*kernel[8];
				ans[6935]<=tmp[6834]*kernel[0]+tmp[6835]*kernel[1]+tmp[6836]*kernel[2]+tmp[6934]*kernel[3]+tmp[6935]*kernel[4]+tmp[6936]*kernel[5]+tmp[7034]*kernel[6]+tmp[7035]*kernel[7]+tmp[7036]*kernel[8];
				ans[6936]<=tmp[6835]*kernel[0]+tmp[6836]*kernel[1]+tmp[6837]*kernel[2]+tmp[6935]*kernel[3]+tmp[6936]*kernel[4]+tmp[6937]*kernel[5]+tmp[7035]*kernel[6]+tmp[7036]*kernel[7]+tmp[7037]*kernel[8];
				ans[6937]<=tmp[6836]*kernel[0]+tmp[6837]*kernel[1]+tmp[6838]*kernel[2]+tmp[6936]*kernel[3]+tmp[6937]*kernel[4]+tmp[6938]*kernel[5]+tmp[7036]*kernel[6]+tmp[7037]*kernel[7]+tmp[7038]*kernel[8];
				ans[6938]<=tmp[6837]*kernel[0]+tmp[6838]*kernel[1]+tmp[6839]*kernel[2]+tmp[6937]*kernel[3]+tmp[6938]*kernel[4]+tmp[6939]*kernel[5]+tmp[7037]*kernel[6]+tmp[7038]*kernel[7]+tmp[7039]*kernel[8];
				ans[6939]<=tmp[6838]*kernel[0]+tmp[6839]*kernel[1]+tmp[6840]*kernel[2]+tmp[6938]*kernel[3]+tmp[6939]*kernel[4]+tmp[6940]*kernel[5]+tmp[7038]*kernel[6]+tmp[7039]*kernel[7]+tmp[7040]*kernel[8];
				ans[6940]<=tmp[6839]*kernel[0]+tmp[6840]*kernel[1]+tmp[6841]*kernel[2]+tmp[6939]*kernel[3]+tmp[6940]*kernel[4]+tmp[6941]*kernel[5]+tmp[7039]*kernel[6]+tmp[7040]*kernel[7]+tmp[7041]*kernel[8];
				ans[6941]<=tmp[6840]*kernel[0]+tmp[6841]*kernel[1]+tmp[6842]*kernel[2]+tmp[6940]*kernel[3]+tmp[6941]*kernel[4]+tmp[6942]*kernel[5]+tmp[7040]*kernel[6]+tmp[7041]*kernel[7]+tmp[7042]*kernel[8];
				ans[6942]<=tmp[6841]*kernel[0]+tmp[6842]*kernel[1]+tmp[6843]*kernel[2]+tmp[6941]*kernel[3]+tmp[6942]*kernel[4]+tmp[6943]*kernel[5]+tmp[7041]*kernel[6]+tmp[7042]*kernel[7]+tmp[7043]*kernel[8];
				ans[6943]<=tmp[6842]*kernel[0]+tmp[6843]*kernel[1]+tmp[6844]*kernel[2]+tmp[6942]*kernel[3]+tmp[6943]*kernel[4]+tmp[6944]*kernel[5]+tmp[7042]*kernel[6]+tmp[7043]*kernel[7]+tmp[7044]*kernel[8];
				ans[6944]<=tmp[6843]*kernel[0]+tmp[6844]*kernel[1]+tmp[6845]*kernel[2]+tmp[6943]*kernel[3]+tmp[6944]*kernel[4]+tmp[6945]*kernel[5]+tmp[7043]*kernel[6]+tmp[7044]*kernel[7]+tmp[7045]*kernel[8];
				ans[6945]<=tmp[6844]*kernel[0]+tmp[6845]*kernel[1]+tmp[6846]*kernel[2]+tmp[6944]*kernel[3]+tmp[6945]*kernel[4]+tmp[6946]*kernel[5]+tmp[7044]*kernel[6]+tmp[7045]*kernel[7]+tmp[7046]*kernel[8];
				ans[6946]<=tmp[6845]*kernel[0]+tmp[6846]*kernel[1]+tmp[6847]*kernel[2]+tmp[6945]*kernel[3]+tmp[6946]*kernel[4]+tmp[6947]*kernel[5]+tmp[7045]*kernel[6]+tmp[7046]*kernel[7]+tmp[7047]*kernel[8];
				ans[6947]<=tmp[6846]*kernel[0]+tmp[6847]*kernel[1]+tmp[6848]*kernel[2]+tmp[6946]*kernel[3]+tmp[6947]*kernel[4]+tmp[6948]*kernel[5]+tmp[7046]*kernel[6]+tmp[7047]*kernel[7]+tmp[7048]*kernel[8];
				ans[6948]<=tmp[6847]*kernel[0]+tmp[6848]*kernel[1]+tmp[6849]*kernel[2]+tmp[6947]*kernel[3]+tmp[6948]*kernel[4]+tmp[6949]*kernel[5]+tmp[7047]*kernel[6]+tmp[7048]*kernel[7]+tmp[7049]*kernel[8];
				ans[6949]<=tmp[6848]*kernel[0]+tmp[6849]*kernel[1]+tmp[6850]*kernel[2]+tmp[6948]*kernel[3]+tmp[6949]*kernel[4]+tmp[6950]*kernel[5]+tmp[7048]*kernel[6]+tmp[7049]*kernel[7]+tmp[7050]*kernel[8];
				ans[6950]<=tmp[6849]*kernel[0]+tmp[6850]*kernel[1]+tmp[6851]*kernel[2]+tmp[6949]*kernel[3]+tmp[6950]*kernel[4]+tmp[6951]*kernel[5]+tmp[7049]*kernel[6]+tmp[7050]*kernel[7]+tmp[7051]*kernel[8];
				ans[6951]<=tmp[6850]*kernel[0]+tmp[6851]*kernel[1]+tmp[6852]*kernel[2]+tmp[6950]*kernel[3]+tmp[6951]*kernel[4]+tmp[6952]*kernel[5]+tmp[7050]*kernel[6]+tmp[7051]*kernel[7]+tmp[7052]*kernel[8];
				ans[6952]<=tmp[6851]*kernel[0]+tmp[6852]*kernel[1]+tmp[6853]*kernel[2]+tmp[6951]*kernel[3]+tmp[6952]*kernel[4]+tmp[6953]*kernel[5]+tmp[7051]*kernel[6]+tmp[7052]*kernel[7]+tmp[7053]*kernel[8];
				ans[6953]<=tmp[6852]*kernel[0]+tmp[6853]*kernel[1]+tmp[6854]*kernel[2]+tmp[6952]*kernel[3]+tmp[6953]*kernel[4]+tmp[6954]*kernel[5]+tmp[7052]*kernel[6]+tmp[7053]*kernel[7]+tmp[7054]*kernel[8];
				ans[6954]<=tmp[6853]*kernel[0]+tmp[6854]*kernel[1]+tmp[6855]*kernel[2]+tmp[6953]*kernel[3]+tmp[6954]*kernel[4]+tmp[6955]*kernel[5]+tmp[7053]*kernel[6]+tmp[7054]*kernel[7]+tmp[7055]*kernel[8];
				ans[6955]<=tmp[6854]*kernel[0]+tmp[6855]*kernel[1]+tmp[6856]*kernel[2]+tmp[6954]*kernel[3]+tmp[6955]*kernel[4]+tmp[6956]*kernel[5]+tmp[7054]*kernel[6]+tmp[7055]*kernel[7]+tmp[7056]*kernel[8];
				ans[6956]<=tmp[6855]*kernel[0]+tmp[6856]*kernel[1]+tmp[6857]*kernel[2]+tmp[6955]*kernel[3]+tmp[6956]*kernel[4]+tmp[6957]*kernel[5]+tmp[7055]*kernel[6]+tmp[7056]*kernel[7]+tmp[7057]*kernel[8];
				ans[6957]<=tmp[6856]*kernel[0]+tmp[6857]*kernel[1]+tmp[6858]*kernel[2]+tmp[6956]*kernel[3]+tmp[6957]*kernel[4]+tmp[6958]*kernel[5]+tmp[7056]*kernel[6]+tmp[7057]*kernel[7]+tmp[7058]*kernel[8];
				ans[6958]<=tmp[6857]*kernel[0]+tmp[6858]*kernel[1]+tmp[6859]*kernel[2]+tmp[6957]*kernel[3]+tmp[6958]*kernel[4]+tmp[6959]*kernel[5]+tmp[7057]*kernel[6]+tmp[7058]*kernel[7]+tmp[7059]*kernel[8];
				ans[6959]<=tmp[6858]*kernel[0]+tmp[6859]*kernel[1]+tmp[6860]*kernel[2]+tmp[6958]*kernel[3]+tmp[6959]*kernel[4]+tmp[6960]*kernel[5]+tmp[7058]*kernel[6]+tmp[7059]*kernel[7]+tmp[7060]*kernel[8];
				ans[6960]<=tmp[6859]*kernel[0]+tmp[6860]*kernel[1]+tmp[6861]*kernel[2]+tmp[6959]*kernel[3]+tmp[6960]*kernel[4]+tmp[6961]*kernel[5]+tmp[7059]*kernel[6]+tmp[7060]*kernel[7]+tmp[7061]*kernel[8];
				ans[6961]<=tmp[6860]*kernel[0]+tmp[6861]*kernel[1]+tmp[6862]*kernel[2]+tmp[6960]*kernel[3]+tmp[6961]*kernel[4]+tmp[6962]*kernel[5]+tmp[7060]*kernel[6]+tmp[7061]*kernel[7]+tmp[7062]*kernel[8];
				ans[6962]<=tmp[6861]*kernel[0]+tmp[6862]*kernel[1]+tmp[6863]*kernel[2]+tmp[6961]*kernel[3]+tmp[6962]*kernel[4]+tmp[6963]*kernel[5]+tmp[7061]*kernel[6]+tmp[7062]*kernel[7]+tmp[7063]*kernel[8];
				ans[6963]<=tmp[6862]*kernel[0]+tmp[6863]*kernel[1]+tmp[6864]*kernel[2]+tmp[6962]*kernel[3]+tmp[6963]*kernel[4]+tmp[6964]*kernel[5]+tmp[7062]*kernel[6]+tmp[7063]*kernel[7]+tmp[7064]*kernel[8];
				ans[6964]<=tmp[6863]*kernel[0]+tmp[6864]*kernel[1]+tmp[6865]*kernel[2]+tmp[6963]*kernel[3]+tmp[6964]*kernel[4]+tmp[6965]*kernel[5]+tmp[7063]*kernel[6]+tmp[7064]*kernel[7]+tmp[7065]*kernel[8];
				ans[6965]<=tmp[6864]*kernel[0]+tmp[6865]*kernel[1]+tmp[6866]*kernel[2]+tmp[6964]*kernel[3]+tmp[6965]*kernel[4]+tmp[6966]*kernel[5]+tmp[7064]*kernel[6]+tmp[7065]*kernel[7]+tmp[7066]*kernel[8];
				ans[6966]<=tmp[6865]*kernel[0]+tmp[6866]*kernel[1]+tmp[6867]*kernel[2]+tmp[6965]*kernel[3]+tmp[6966]*kernel[4]+tmp[6967]*kernel[5]+tmp[7065]*kernel[6]+tmp[7066]*kernel[7]+tmp[7067]*kernel[8];
				ans[6967]<=tmp[6866]*kernel[0]+tmp[6867]*kernel[1]+tmp[6868]*kernel[2]+tmp[6966]*kernel[3]+tmp[6967]*kernel[4]+tmp[6968]*kernel[5]+tmp[7066]*kernel[6]+tmp[7067]*kernel[7]+tmp[7068]*kernel[8];
				ans[6968]<=tmp[6867]*kernel[0]+tmp[6868]*kernel[1]+tmp[6869]*kernel[2]+tmp[6967]*kernel[3]+tmp[6968]*kernel[4]+tmp[6969]*kernel[5]+tmp[7067]*kernel[6]+tmp[7068]*kernel[7]+tmp[7069]*kernel[8];
				ans[6969]<=tmp[6868]*kernel[0]+tmp[6869]*kernel[1]+tmp[6870]*kernel[2]+tmp[6968]*kernel[3]+tmp[6969]*kernel[4]+tmp[6970]*kernel[5]+tmp[7068]*kernel[6]+tmp[7069]*kernel[7]+tmp[7070]*kernel[8];
				ans[6970]<=tmp[6869]*kernel[0]+tmp[6870]*kernel[1]+tmp[6871]*kernel[2]+tmp[6969]*kernel[3]+tmp[6970]*kernel[4]+tmp[6971]*kernel[5]+tmp[7069]*kernel[6]+tmp[7070]*kernel[7]+tmp[7071]*kernel[8];
				ans[6971]<=tmp[6870]*kernel[0]+tmp[6871]*kernel[1]+tmp[6872]*kernel[2]+tmp[6970]*kernel[3]+tmp[6971]*kernel[4]+tmp[6972]*kernel[5]+tmp[7070]*kernel[6]+tmp[7071]*kernel[7]+tmp[7072]*kernel[8];
				ans[6972]<=tmp[6871]*kernel[0]+tmp[6872]*kernel[1]+tmp[6873]*kernel[2]+tmp[6971]*kernel[3]+tmp[6972]*kernel[4]+tmp[6973]*kernel[5]+tmp[7071]*kernel[6]+tmp[7072]*kernel[7]+tmp[7073]*kernel[8];
				ans[6973]<=tmp[6872]*kernel[0]+tmp[6873]*kernel[1]+tmp[6874]*kernel[2]+tmp[6972]*kernel[3]+tmp[6973]*kernel[4]+tmp[6974]*kernel[5]+tmp[7072]*kernel[6]+tmp[7073]*kernel[7]+tmp[7074]*kernel[8];
				ans[6974]<=tmp[6873]*kernel[0]+tmp[6874]*kernel[1]+tmp[6875]*kernel[2]+tmp[6973]*kernel[3]+tmp[6974]*kernel[4]+tmp[6975]*kernel[5]+tmp[7073]*kernel[6]+tmp[7074]*kernel[7]+tmp[7075]*kernel[8];
				ans[6975]<=tmp[6874]*kernel[0]+tmp[6875]*kernel[1]+tmp[6876]*kernel[2]+tmp[6974]*kernel[3]+tmp[6975]*kernel[4]+tmp[6976]*kernel[5]+tmp[7074]*kernel[6]+tmp[7075]*kernel[7]+tmp[7076]*kernel[8];
				ans[6976]<=tmp[6875]*kernel[0]+tmp[6876]*kernel[1]+tmp[6877]*kernel[2]+tmp[6975]*kernel[3]+tmp[6976]*kernel[4]+tmp[6977]*kernel[5]+tmp[7075]*kernel[6]+tmp[7076]*kernel[7]+tmp[7077]*kernel[8];
				ans[6977]<=tmp[6876]*kernel[0]+tmp[6877]*kernel[1]+tmp[6878]*kernel[2]+tmp[6976]*kernel[3]+tmp[6977]*kernel[4]+tmp[6978]*kernel[5]+tmp[7076]*kernel[6]+tmp[7077]*kernel[7]+tmp[7078]*kernel[8];
				ans[6978]<=tmp[6877]*kernel[0]+tmp[6878]*kernel[1]+tmp[6879]*kernel[2]+tmp[6977]*kernel[3]+tmp[6978]*kernel[4]+tmp[6979]*kernel[5]+tmp[7077]*kernel[6]+tmp[7078]*kernel[7]+tmp[7079]*kernel[8];
				ans[6979]<=tmp[6878]*kernel[0]+tmp[6879]*kernel[1]+tmp[6880]*kernel[2]+tmp[6978]*kernel[3]+tmp[6979]*kernel[4]+tmp[6980]*kernel[5]+tmp[7078]*kernel[6]+tmp[7079]*kernel[7]+tmp[7080]*kernel[8];
				ans[6980]<=tmp[6879]*kernel[0]+tmp[6880]*kernel[1]+tmp[6881]*kernel[2]+tmp[6979]*kernel[3]+tmp[6980]*kernel[4]+tmp[6981]*kernel[5]+tmp[7079]*kernel[6]+tmp[7080]*kernel[7]+tmp[7081]*kernel[8];
				ans[6981]<=tmp[6880]*kernel[0]+tmp[6881]*kernel[1]+tmp[6882]*kernel[2]+tmp[6980]*kernel[3]+tmp[6981]*kernel[4]+tmp[6982]*kernel[5]+tmp[7080]*kernel[6]+tmp[7081]*kernel[7]+tmp[7082]*kernel[8];
				ans[6982]<=tmp[6881]*kernel[0]+tmp[6882]*kernel[1]+tmp[6883]*kernel[2]+tmp[6981]*kernel[3]+tmp[6982]*kernel[4]+tmp[6983]*kernel[5]+tmp[7081]*kernel[6]+tmp[7082]*kernel[7]+tmp[7083]*kernel[8];
				ans[6983]<=tmp[6882]*kernel[0]+tmp[6883]*kernel[1]+tmp[6884]*kernel[2]+tmp[6982]*kernel[3]+tmp[6983]*kernel[4]+tmp[6984]*kernel[5]+tmp[7082]*kernel[6]+tmp[7083]*kernel[7]+tmp[7084]*kernel[8];
				ans[6984]<=tmp[6883]*kernel[0]+tmp[6884]*kernel[1]+tmp[6885]*kernel[2]+tmp[6983]*kernel[3]+tmp[6984]*kernel[4]+tmp[6985]*kernel[5]+tmp[7083]*kernel[6]+tmp[7084]*kernel[7]+tmp[7085]*kernel[8];
				ans[6985]<=tmp[6884]*kernel[0]+tmp[6885]*kernel[1]+tmp[6886]*kernel[2]+tmp[6984]*kernel[3]+tmp[6985]*kernel[4]+tmp[6986]*kernel[5]+tmp[7084]*kernel[6]+tmp[7085]*kernel[7]+tmp[7086]*kernel[8];
				ans[6986]<=tmp[6885]*kernel[0]+tmp[6886]*kernel[1]+tmp[6887]*kernel[2]+tmp[6985]*kernel[3]+tmp[6986]*kernel[4]+tmp[6987]*kernel[5]+tmp[7085]*kernel[6]+tmp[7086]*kernel[7]+tmp[7087]*kernel[8];
				ans[6987]<=tmp[6886]*kernel[0]+tmp[6887]*kernel[1]+tmp[6888]*kernel[2]+tmp[6986]*kernel[3]+tmp[6987]*kernel[4]+tmp[6988]*kernel[5]+tmp[7086]*kernel[6]+tmp[7087]*kernel[7]+tmp[7088]*kernel[8];
				ans[6988]<=tmp[6887]*kernel[0]+tmp[6888]*kernel[1]+tmp[6889]*kernel[2]+tmp[6987]*kernel[3]+tmp[6988]*kernel[4]+tmp[6989]*kernel[5]+tmp[7087]*kernel[6]+tmp[7088]*kernel[7]+tmp[7089]*kernel[8];
				ans[6989]<=tmp[6888]*kernel[0]+tmp[6889]*kernel[1]+tmp[6890]*kernel[2]+tmp[6988]*kernel[3]+tmp[6989]*kernel[4]+tmp[6990]*kernel[5]+tmp[7088]*kernel[6]+tmp[7089]*kernel[7]+tmp[7090]*kernel[8];
				ans[6990]<=tmp[6889]*kernel[0]+tmp[6890]*kernel[1]+tmp[6891]*kernel[2]+tmp[6989]*kernel[3]+tmp[6990]*kernel[4]+tmp[6991]*kernel[5]+tmp[7089]*kernel[6]+tmp[7090]*kernel[7]+tmp[7091]*kernel[8];
				ans[6991]<=tmp[6890]*kernel[0]+tmp[6891]*kernel[1]+tmp[6892]*kernel[2]+tmp[6990]*kernel[3]+tmp[6991]*kernel[4]+tmp[6992]*kernel[5]+tmp[7090]*kernel[6]+tmp[7091]*kernel[7]+tmp[7092]*kernel[8];
				ans[6992]<=tmp[6891]*kernel[0]+tmp[6892]*kernel[1]+tmp[6893]*kernel[2]+tmp[6991]*kernel[3]+tmp[6992]*kernel[4]+tmp[6993]*kernel[5]+tmp[7091]*kernel[6]+tmp[7092]*kernel[7]+tmp[7093]*kernel[8];
				ans[6993]<=tmp[6892]*kernel[0]+tmp[6893]*kernel[1]+tmp[6894]*kernel[2]+tmp[6992]*kernel[3]+tmp[6993]*kernel[4]+tmp[6994]*kernel[5]+tmp[7092]*kernel[6]+tmp[7093]*kernel[7]+tmp[7094]*kernel[8];
				ans[6994]<=tmp[6893]*kernel[0]+tmp[6894]*kernel[1]+tmp[6895]*kernel[2]+tmp[6993]*kernel[3]+tmp[6994]*kernel[4]+tmp[6995]*kernel[5]+tmp[7093]*kernel[6]+tmp[7094]*kernel[7]+tmp[7095]*kernel[8];
				ans[6995]<=tmp[6894]*kernel[0]+tmp[6895]*kernel[1]+tmp[6896]*kernel[2]+tmp[6994]*kernel[3]+tmp[6995]*kernel[4]+tmp[6996]*kernel[5]+tmp[7094]*kernel[6]+tmp[7095]*kernel[7]+tmp[7096]*kernel[8];
				ans[6996]<=tmp[6895]*kernel[0]+tmp[6896]*kernel[1]+tmp[6897]*kernel[2]+tmp[6995]*kernel[3]+tmp[6996]*kernel[4]+tmp[6997]*kernel[5]+tmp[7095]*kernel[6]+tmp[7096]*kernel[7]+tmp[7097]*kernel[8];
				ans[6997]<=tmp[6896]*kernel[0]+tmp[6897]*kernel[1]+tmp[6898]*kernel[2]+tmp[6996]*kernel[3]+tmp[6997]*kernel[4]+tmp[6998]*kernel[5]+tmp[7096]*kernel[6]+tmp[7097]*kernel[7]+tmp[7098]*kernel[8];
				ans[6998]<=tmp[6897]*kernel[0]+tmp[6898]*kernel[1]+tmp[6899]*kernel[2]+tmp[6997]*kernel[3]+tmp[6998]*kernel[4]+tmp[6999]*kernel[5]+tmp[7097]*kernel[6]+tmp[7098]*kernel[7]+tmp[7099]*kernel[8];
				ans[6999]<=tmp[6898]*kernel[0]+tmp[6899]*kernel[1]+tmp[6998]*kernel[3]+tmp[6999]*kernel[4]+tmp[7098]*kernel[6]+tmp[7099]*kernel[7];
				ans[7000]<=tmp[6900]*kernel[1]+tmp[6901]*kernel[2]+tmp[7000]*kernel[4]+tmp[7001]*kernel[5]+tmp[7100]*kernel[7]+tmp[7101]*kernel[8];
				ans[7001]<=tmp[6900]*kernel[0]+tmp[6901]*kernel[1]+tmp[6902]*kernel[2]+tmp[7000]*kernel[3]+tmp[7001]*kernel[4]+tmp[7002]*kernel[5]+tmp[7100]*kernel[6]+tmp[7101]*kernel[7]+tmp[7102]*kernel[8];
				ans[7002]<=tmp[6901]*kernel[0]+tmp[6902]*kernel[1]+tmp[6903]*kernel[2]+tmp[7001]*kernel[3]+tmp[7002]*kernel[4]+tmp[7003]*kernel[5]+tmp[7101]*kernel[6]+tmp[7102]*kernel[7]+tmp[7103]*kernel[8];
				ans[7003]<=tmp[6902]*kernel[0]+tmp[6903]*kernel[1]+tmp[6904]*kernel[2]+tmp[7002]*kernel[3]+tmp[7003]*kernel[4]+tmp[7004]*kernel[5]+tmp[7102]*kernel[6]+tmp[7103]*kernel[7]+tmp[7104]*kernel[8];
				ans[7004]<=tmp[6903]*kernel[0]+tmp[6904]*kernel[1]+tmp[6905]*kernel[2]+tmp[7003]*kernel[3]+tmp[7004]*kernel[4]+tmp[7005]*kernel[5]+tmp[7103]*kernel[6]+tmp[7104]*kernel[7]+tmp[7105]*kernel[8];
				ans[7005]<=tmp[6904]*kernel[0]+tmp[6905]*kernel[1]+tmp[6906]*kernel[2]+tmp[7004]*kernel[3]+tmp[7005]*kernel[4]+tmp[7006]*kernel[5]+tmp[7104]*kernel[6]+tmp[7105]*kernel[7]+tmp[7106]*kernel[8];
				ans[7006]<=tmp[6905]*kernel[0]+tmp[6906]*kernel[1]+tmp[6907]*kernel[2]+tmp[7005]*kernel[3]+tmp[7006]*kernel[4]+tmp[7007]*kernel[5]+tmp[7105]*kernel[6]+tmp[7106]*kernel[7]+tmp[7107]*kernel[8];
				ans[7007]<=tmp[6906]*kernel[0]+tmp[6907]*kernel[1]+tmp[6908]*kernel[2]+tmp[7006]*kernel[3]+tmp[7007]*kernel[4]+tmp[7008]*kernel[5]+tmp[7106]*kernel[6]+tmp[7107]*kernel[7]+tmp[7108]*kernel[8];
				ans[7008]<=tmp[6907]*kernel[0]+tmp[6908]*kernel[1]+tmp[6909]*kernel[2]+tmp[7007]*kernel[3]+tmp[7008]*kernel[4]+tmp[7009]*kernel[5]+tmp[7107]*kernel[6]+tmp[7108]*kernel[7]+tmp[7109]*kernel[8];
				ans[7009]<=tmp[6908]*kernel[0]+tmp[6909]*kernel[1]+tmp[6910]*kernel[2]+tmp[7008]*kernel[3]+tmp[7009]*kernel[4]+tmp[7010]*kernel[5]+tmp[7108]*kernel[6]+tmp[7109]*kernel[7]+tmp[7110]*kernel[8];
				ans[7010]<=tmp[6909]*kernel[0]+tmp[6910]*kernel[1]+tmp[6911]*kernel[2]+tmp[7009]*kernel[3]+tmp[7010]*kernel[4]+tmp[7011]*kernel[5]+tmp[7109]*kernel[6]+tmp[7110]*kernel[7]+tmp[7111]*kernel[8];
				ans[7011]<=tmp[6910]*kernel[0]+tmp[6911]*kernel[1]+tmp[6912]*kernel[2]+tmp[7010]*kernel[3]+tmp[7011]*kernel[4]+tmp[7012]*kernel[5]+tmp[7110]*kernel[6]+tmp[7111]*kernel[7]+tmp[7112]*kernel[8];
				ans[7012]<=tmp[6911]*kernel[0]+tmp[6912]*kernel[1]+tmp[6913]*kernel[2]+tmp[7011]*kernel[3]+tmp[7012]*kernel[4]+tmp[7013]*kernel[5]+tmp[7111]*kernel[6]+tmp[7112]*kernel[7]+tmp[7113]*kernel[8];
				ans[7013]<=tmp[6912]*kernel[0]+tmp[6913]*kernel[1]+tmp[6914]*kernel[2]+tmp[7012]*kernel[3]+tmp[7013]*kernel[4]+tmp[7014]*kernel[5]+tmp[7112]*kernel[6]+tmp[7113]*kernel[7]+tmp[7114]*kernel[8];
				ans[7014]<=tmp[6913]*kernel[0]+tmp[6914]*kernel[1]+tmp[6915]*kernel[2]+tmp[7013]*kernel[3]+tmp[7014]*kernel[4]+tmp[7015]*kernel[5]+tmp[7113]*kernel[6]+tmp[7114]*kernel[7]+tmp[7115]*kernel[8];
				ans[7015]<=tmp[6914]*kernel[0]+tmp[6915]*kernel[1]+tmp[6916]*kernel[2]+tmp[7014]*kernel[3]+tmp[7015]*kernel[4]+tmp[7016]*kernel[5]+tmp[7114]*kernel[6]+tmp[7115]*kernel[7]+tmp[7116]*kernel[8];
				ans[7016]<=tmp[6915]*kernel[0]+tmp[6916]*kernel[1]+tmp[6917]*kernel[2]+tmp[7015]*kernel[3]+tmp[7016]*kernel[4]+tmp[7017]*kernel[5]+tmp[7115]*kernel[6]+tmp[7116]*kernel[7]+tmp[7117]*kernel[8];
				ans[7017]<=tmp[6916]*kernel[0]+tmp[6917]*kernel[1]+tmp[6918]*kernel[2]+tmp[7016]*kernel[3]+tmp[7017]*kernel[4]+tmp[7018]*kernel[5]+tmp[7116]*kernel[6]+tmp[7117]*kernel[7]+tmp[7118]*kernel[8];
				ans[7018]<=tmp[6917]*kernel[0]+tmp[6918]*kernel[1]+tmp[6919]*kernel[2]+tmp[7017]*kernel[3]+tmp[7018]*kernel[4]+tmp[7019]*kernel[5]+tmp[7117]*kernel[6]+tmp[7118]*kernel[7]+tmp[7119]*kernel[8];
				ans[7019]<=tmp[6918]*kernel[0]+tmp[6919]*kernel[1]+tmp[6920]*kernel[2]+tmp[7018]*kernel[3]+tmp[7019]*kernel[4]+tmp[7020]*kernel[5]+tmp[7118]*kernel[6]+tmp[7119]*kernel[7]+tmp[7120]*kernel[8];
				ans[7020]<=tmp[6919]*kernel[0]+tmp[6920]*kernel[1]+tmp[6921]*kernel[2]+tmp[7019]*kernel[3]+tmp[7020]*kernel[4]+tmp[7021]*kernel[5]+tmp[7119]*kernel[6]+tmp[7120]*kernel[7]+tmp[7121]*kernel[8];
				ans[7021]<=tmp[6920]*kernel[0]+tmp[6921]*kernel[1]+tmp[6922]*kernel[2]+tmp[7020]*kernel[3]+tmp[7021]*kernel[4]+tmp[7022]*kernel[5]+tmp[7120]*kernel[6]+tmp[7121]*kernel[7]+tmp[7122]*kernel[8];
				ans[7022]<=tmp[6921]*kernel[0]+tmp[6922]*kernel[1]+tmp[6923]*kernel[2]+tmp[7021]*kernel[3]+tmp[7022]*kernel[4]+tmp[7023]*kernel[5]+tmp[7121]*kernel[6]+tmp[7122]*kernel[7]+tmp[7123]*kernel[8];
				ans[7023]<=tmp[6922]*kernel[0]+tmp[6923]*kernel[1]+tmp[6924]*kernel[2]+tmp[7022]*kernel[3]+tmp[7023]*kernel[4]+tmp[7024]*kernel[5]+tmp[7122]*kernel[6]+tmp[7123]*kernel[7]+tmp[7124]*kernel[8];
				ans[7024]<=tmp[6923]*kernel[0]+tmp[6924]*kernel[1]+tmp[6925]*kernel[2]+tmp[7023]*kernel[3]+tmp[7024]*kernel[4]+tmp[7025]*kernel[5]+tmp[7123]*kernel[6]+tmp[7124]*kernel[7]+tmp[7125]*kernel[8];
				ans[7025]<=tmp[6924]*kernel[0]+tmp[6925]*kernel[1]+tmp[6926]*kernel[2]+tmp[7024]*kernel[3]+tmp[7025]*kernel[4]+tmp[7026]*kernel[5]+tmp[7124]*kernel[6]+tmp[7125]*kernel[7]+tmp[7126]*kernel[8];
				ans[7026]<=tmp[6925]*kernel[0]+tmp[6926]*kernel[1]+tmp[6927]*kernel[2]+tmp[7025]*kernel[3]+tmp[7026]*kernel[4]+tmp[7027]*kernel[5]+tmp[7125]*kernel[6]+tmp[7126]*kernel[7]+tmp[7127]*kernel[8];
				ans[7027]<=tmp[6926]*kernel[0]+tmp[6927]*kernel[1]+tmp[6928]*kernel[2]+tmp[7026]*kernel[3]+tmp[7027]*kernel[4]+tmp[7028]*kernel[5]+tmp[7126]*kernel[6]+tmp[7127]*kernel[7]+tmp[7128]*kernel[8];
				ans[7028]<=tmp[6927]*kernel[0]+tmp[6928]*kernel[1]+tmp[6929]*kernel[2]+tmp[7027]*kernel[3]+tmp[7028]*kernel[4]+tmp[7029]*kernel[5]+tmp[7127]*kernel[6]+tmp[7128]*kernel[7]+tmp[7129]*kernel[8];
				ans[7029]<=tmp[6928]*kernel[0]+tmp[6929]*kernel[1]+tmp[6930]*kernel[2]+tmp[7028]*kernel[3]+tmp[7029]*kernel[4]+tmp[7030]*kernel[5]+tmp[7128]*kernel[6]+tmp[7129]*kernel[7]+tmp[7130]*kernel[8];
				ans[7030]<=tmp[6929]*kernel[0]+tmp[6930]*kernel[1]+tmp[6931]*kernel[2]+tmp[7029]*kernel[3]+tmp[7030]*kernel[4]+tmp[7031]*kernel[5]+tmp[7129]*kernel[6]+tmp[7130]*kernel[7]+tmp[7131]*kernel[8];
				ans[7031]<=tmp[6930]*kernel[0]+tmp[6931]*kernel[1]+tmp[6932]*kernel[2]+tmp[7030]*kernel[3]+tmp[7031]*kernel[4]+tmp[7032]*kernel[5]+tmp[7130]*kernel[6]+tmp[7131]*kernel[7]+tmp[7132]*kernel[8];
				ans[7032]<=tmp[6931]*kernel[0]+tmp[6932]*kernel[1]+tmp[6933]*kernel[2]+tmp[7031]*kernel[3]+tmp[7032]*kernel[4]+tmp[7033]*kernel[5]+tmp[7131]*kernel[6]+tmp[7132]*kernel[7]+tmp[7133]*kernel[8];
				ans[7033]<=tmp[6932]*kernel[0]+tmp[6933]*kernel[1]+tmp[6934]*kernel[2]+tmp[7032]*kernel[3]+tmp[7033]*kernel[4]+tmp[7034]*kernel[5]+tmp[7132]*kernel[6]+tmp[7133]*kernel[7]+tmp[7134]*kernel[8];
				ans[7034]<=tmp[6933]*kernel[0]+tmp[6934]*kernel[1]+tmp[6935]*kernel[2]+tmp[7033]*kernel[3]+tmp[7034]*kernel[4]+tmp[7035]*kernel[5]+tmp[7133]*kernel[6]+tmp[7134]*kernel[7]+tmp[7135]*kernel[8];
				ans[7035]<=tmp[6934]*kernel[0]+tmp[6935]*kernel[1]+tmp[6936]*kernel[2]+tmp[7034]*kernel[3]+tmp[7035]*kernel[4]+tmp[7036]*kernel[5]+tmp[7134]*kernel[6]+tmp[7135]*kernel[7]+tmp[7136]*kernel[8];
				ans[7036]<=tmp[6935]*kernel[0]+tmp[6936]*kernel[1]+tmp[6937]*kernel[2]+tmp[7035]*kernel[3]+tmp[7036]*kernel[4]+tmp[7037]*kernel[5]+tmp[7135]*kernel[6]+tmp[7136]*kernel[7]+tmp[7137]*kernel[8];
				ans[7037]<=tmp[6936]*kernel[0]+tmp[6937]*kernel[1]+tmp[6938]*kernel[2]+tmp[7036]*kernel[3]+tmp[7037]*kernel[4]+tmp[7038]*kernel[5]+tmp[7136]*kernel[6]+tmp[7137]*kernel[7]+tmp[7138]*kernel[8];
				ans[7038]<=tmp[6937]*kernel[0]+tmp[6938]*kernel[1]+tmp[6939]*kernel[2]+tmp[7037]*kernel[3]+tmp[7038]*kernel[4]+tmp[7039]*kernel[5]+tmp[7137]*kernel[6]+tmp[7138]*kernel[7]+tmp[7139]*kernel[8];
				ans[7039]<=tmp[6938]*kernel[0]+tmp[6939]*kernel[1]+tmp[6940]*kernel[2]+tmp[7038]*kernel[3]+tmp[7039]*kernel[4]+tmp[7040]*kernel[5]+tmp[7138]*kernel[6]+tmp[7139]*kernel[7]+tmp[7140]*kernel[8];
				ans[7040]<=tmp[6939]*kernel[0]+tmp[6940]*kernel[1]+tmp[6941]*kernel[2]+tmp[7039]*kernel[3]+tmp[7040]*kernel[4]+tmp[7041]*kernel[5]+tmp[7139]*kernel[6]+tmp[7140]*kernel[7]+tmp[7141]*kernel[8];
				ans[7041]<=tmp[6940]*kernel[0]+tmp[6941]*kernel[1]+tmp[6942]*kernel[2]+tmp[7040]*kernel[3]+tmp[7041]*kernel[4]+tmp[7042]*kernel[5]+tmp[7140]*kernel[6]+tmp[7141]*kernel[7]+tmp[7142]*kernel[8];
				ans[7042]<=tmp[6941]*kernel[0]+tmp[6942]*kernel[1]+tmp[6943]*kernel[2]+tmp[7041]*kernel[3]+tmp[7042]*kernel[4]+tmp[7043]*kernel[5]+tmp[7141]*kernel[6]+tmp[7142]*kernel[7]+tmp[7143]*kernel[8];
				ans[7043]<=tmp[6942]*kernel[0]+tmp[6943]*kernel[1]+tmp[6944]*kernel[2]+tmp[7042]*kernel[3]+tmp[7043]*kernel[4]+tmp[7044]*kernel[5]+tmp[7142]*kernel[6]+tmp[7143]*kernel[7]+tmp[7144]*kernel[8];
				ans[7044]<=tmp[6943]*kernel[0]+tmp[6944]*kernel[1]+tmp[6945]*kernel[2]+tmp[7043]*kernel[3]+tmp[7044]*kernel[4]+tmp[7045]*kernel[5]+tmp[7143]*kernel[6]+tmp[7144]*kernel[7]+tmp[7145]*kernel[8];
				ans[7045]<=tmp[6944]*kernel[0]+tmp[6945]*kernel[1]+tmp[6946]*kernel[2]+tmp[7044]*kernel[3]+tmp[7045]*kernel[4]+tmp[7046]*kernel[5]+tmp[7144]*kernel[6]+tmp[7145]*kernel[7]+tmp[7146]*kernel[8];
				ans[7046]<=tmp[6945]*kernel[0]+tmp[6946]*kernel[1]+tmp[6947]*kernel[2]+tmp[7045]*kernel[3]+tmp[7046]*kernel[4]+tmp[7047]*kernel[5]+tmp[7145]*kernel[6]+tmp[7146]*kernel[7]+tmp[7147]*kernel[8];
				ans[7047]<=tmp[6946]*kernel[0]+tmp[6947]*kernel[1]+tmp[6948]*kernel[2]+tmp[7046]*kernel[3]+tmp[7047]*kernel[4]+tmp[7048]*kernel[5]+tmp[7146]*kernel[6]+tmp[7147]*kernel[7]+tmp[7148]*kernel[8];
				ans[7048]<=tmp[6947]*kernel[0]+tmp[6948]*kernel[1]+tmp[6949]*kernel[2]+tmp[7047]*kernel[3]+tmp[7048]*kernel[4]+tmp[7049]*kernel[5]+tmp[7147]*kernel[6]+tmp[7148]*kernel[7]+tmp[7149]*kernel[8];
				ans[7049]<=tmp[6948]*kernel[0]+tmp[6949]*kernel[1]+tmp[6950]*kernel[2]+tmp[7048]*kernel[3]+tmp[7049]*kernel[4]+tmp[7050]*kernel[5]+tmp[7148]*kernel[6]+tmp[7149]*kernel[7]+tmp[7150]*kernel[8];
				ans[7050]<=tmp[6949]*kernel[0]+tmp[6950]*kernel[1]+tmp[6951]*kernel[2]+tmp[7049]*kernel[3]+tmp[7050]*kernel[4]+tmp[7051]*kernel[5]+tmp[7149]*kernel[6]+tmp[7150]*kernel[7]+tmp[7151]*kernel[8];
				ans[7051]<=tmp[6950]*kernel[0]+tmp[6951]*kernel[1]+tmp[6952]*kernel[2]+tmp[7050]*kernel[3]+tmp[7051]*kernel[4]+tmp[7052]*kernel[5]+tmp[7150]*kernel[6]+tmp[7151]*kernel[7]+tmp[7152]*kernel[8];
				ans[7052]<=tmp[6951]*kernel[0]+tmp[6952]*kernel[1]+tmp[6953]*kernel[2]+tmp[7051]*kernel[3]+tmp[7052]*kernel[4]+tmp[7053]*kernel[5]+tmp[7151]*kernel[6]+tmp[7152]*kernel[7]+tmp[7153]*kernel[8];
				ans[7053]<=tmp[6952]*kernel[0]+tmp[6953]*kernel[1]+tmp[6954]*kernel[2]+tmp[7052]*kernel[3]+tmp[7053]*kernel[4]+tmp[7054]*kernel[5]+tmp[7152]*kernel[6]+tmp[7153]*kernel[7]+tmp[7154]*kernel[8];
				ans[7054]<=tmp[6953]*kernel[0]+tmp[6954]*kernel[1]+tmp[6955]*kernel[2]+tmp[7053]*kernel[3]+tmp[7054]*kernel[4]+tmp[7055]*kernel[5]+tmp[7153]*kernel[6]+tmp[7154]*kernel[7]+tmp[7155]*kernel[8];
				ans[7055]<=tmp[6954]*kernel[0]+tmp[6955]*kernel[1]+tmp[6956]*kernel[2]+tmp[7054]*kernel[3]+tmp[7055]*kernel[4]+tmp[7056]*kernel[5]+tmp[7154]*kernel[6]+tmp[7155]*kernel[7]+tmp[7156]*kernel[8];
				ans[7056]<=tmp[6955]*kernel[0]+tmp[6956]*kernel[1]+tmp[6957]*kernel[2]+tmp[7055]*kernel[3]+tmp[7056]*kernel[4]+tmp[7057]*kernel[5]+tmp[7155]*kernel[6]+tmp[7156]*kernel[7]+tmp[7157]*kernel[8];
				ans[7057]<=tmp[6956]*kernel[0]+tmp[6957]*kernel[1]+tmp[6958]*kernel[2]+tmp[7056]*kernel[3]+tmp[7057]*kernel[4]+tmp[7058]*kernel[5]+tmp[7156]*kernel[6]+tmp[7157]*kernel[7]+tmp[7158]*kernel[8];
				ans[7058]<=tmp[6957]*kernel[0]+tmp[6958]*kernel[1]+tmp[6959]*kernel[2]+tmp[7057]*kernel[3]+tmp[7058]*kernel[4]+tmp[7059]*kernel[5]+tmp[7157]*kernel[6]+tmp[7158]*kernel[7]+tmp[7159]*kernel[8];
				ans[7059]<=tmp[6958]*kernel[0]+tmp[6959]*kernel[1]+tmp[6960]*kernel[2]+tmp[7058]*kernel[3]+tmp[7059]*kernel[4]+tmp[7060]*kernel[5]+tmp[7158]*kernel[6]+tmp[7159]*kernel[7]+tmp[7160]*kernel[8];
				ans[7060]<=tmp[6959]*kernel[0]+tmp[6960]*kernel[1]+tmp[6961]*kernel[2]+tmp[7059]*kernel[3]+tmp[7060]*kernel[4]+tmp[7061]*kernel[5]+tmp[7159]*kernel[6]+tmp[7160]*kernel[7]+tmp[7161]*kernel[8];
				ans[7061]<=tmp[6960]*kernel[0]+tmp[6961]*kernel[1]+tmp[6962]*kernel[2]+tmp[7060]*kernel[3]+tmp[7061]*kernel[4]+tmp[7062]*kernel[5]+tmp[7160]*kernel[6]+tmp[7161]*kernel[7]+tmp[7162]*kernel[8];
				ans[7062]<=tmp[6961]*kernel[0]+tmp[6962]*kernel[1]+tmp[6963]*kernel[2]+tmp[7061]*kernel[3]+tmp[7062]*kernel[4]+tmp[7063]*kernel[5]+tmp[7161]*kernel[6]+tmp[7162]*kernel[7]+tmp[7163]*kernel[8];
				ans[7063]<=tmp[6962]*kernel[0]+tmp[6963]*kernel[1]+tmp[6964]*kernel[2]+tmp[7062]*kernel[3]+tmp[7063]*kernel[4]+tmp[7064]*kernel[5]+tmp[7162]*kernel[6]+tmp[7163]*kernel[7]+tmp[7164]*kernel[8];
				ans[7064]<=tmp[6963]*kernel[0]+tmp[6964]*kernel[1]+tmp[6965]*kernel[2]+tmp[7063]*kernel[3]+tmp[7064]*kernel[4]+tmp[7065]*kernel[5]+tmp[7163]*kernel[6]+tmp[7164]*kernel[7]+tmp[7165]*kernel[8];
				ans[7065]<=tmp[6964]*kernel[0]+tmp[6965]*kernel[1]+tmp[6966]*kernel[2]+tmp[7064]*kernel[3]+tmp[7065]*kernel[4]+tmp[7066]*kernel[5]+tmp[7164]*kernel[6]+tmp[7165]*kernel[7]+tmp[7166]*kernel[8];
				ans[7066]<=tmp[6965]*kernel[0]+tmp[6966]*kernel[1]+tmp[6967]*kernel[2]+tmp[7065]*kernel[3]+tmp[7066]*kernel[4]+tmp[7067]*kernel[5]+tmp[7165]*kernel[6]+tmp[7166]*kernel[7]+tmp[7167]*kernel[8];
				ans[7067]<=tmp[6966]*kernel[0]+tmp[6967]*kernel[1]+tmp[6968]*kernel[2]+tmp[7066]*kernel[3]+tmp[7067]*kernel[4]+tmp[7068]*kernel[5]+tmp[7166]*kernel[6]+tmp[7167]*kernel[7]+tmp[7168]*kernel[8];
				ans[7068]<=tmp[6967]*kernel[0]+tmp[6968]*kernel[1]+tmp[6969]*kernel[2]+tmp[7067]*kernel[3]+tmp[7068]*kernel[4]+tmp[7069]*kernel[5]+tmp[7167]*kernel[6]+tmp[7168]*kernel[7]+tmp[7169]*kernel[8];
				ans[7069]<=tmp[6968]*kernel[0]+tmp[6969]*kernel[1]+tmp[6970]*kernel[2]+tmp[7068]*kernel[3]+tmp[7069]*kernel[4]+tmp[7070]*kernel[5]+tmp[7168]*kernel[6]+tmp[7169]*kernel[7]+tmp[7170]*kernel[8];
				ans[7070]<=tmp[6969]*kernel[0]+tmp[6970]*kernel[1]+tmp[6971]*kernel[2]+tmp[7069]*kernel[3]+tmp[7070]*kernel[4]+tmp[7071]*kernel[5]+tmp[7169]*kernel[6]+tmp[7170]*kernel[7]+tmp[7171]*kernel[8];
				ans[7071]<=tmp[6970]*kernel[0]+tmp[6971]*kernel[1]+tmp[6972]*kernel[2]+tmp[7070]*kernel[3]+tmp[7071]*kernel[4]+tmp[7072]*kernel[5]+tmp[7170]*kernel[6]+tmp[7171]*kernel[7]+tmp[7172]*kernel[8];
				ans[7072]<=tmp[6971]*kernel[0]+tmp[6972]*kernel[1]+tmp[6973]*kernel[2]+tmp[7071]*kernel[3]+tmp[7072]*kernel[4]+tmp[7073]*kernel[5]+tmp[7171]*kernel[6]+tmp[7172]*kernel[7]+tmp[7173]*kernel[8];
				ans[7073]<=tmp[6972]*kernel[0]+tmp[6973]*kernel[1]+tmp[6974]*kernel[2]+tmp[7072]*kernel[3]+tmp[7073]*kernel[4]+tmp[7074]*kernel[5]+tmp[7172]*kernel[6]+tmp[7173]*kernel[7]+tmp[7174]*kernel[8];
				ans[7074]<=tmp[6973]*kernel[0]+tmp[6974]*kernel[1]+tmp[6975]*kernel[2]+tmp[7073]*kernel[3]+tmp[7074]*kernel[4]+tmp[7075]*kernel[5]+tmp[7173]*kernel[6]+tmp[7174]*kernel[7]+tmp[7175]*kernel[8];
				ans[7075]<=tmp[6974]*kernel[0]+tmp[6975]*kernel[1]+tmp[6976]*kernel[2]+tmp[7074]*kernel[3]+tmp[7075]*kernel[4]+tmp[7076]*kernel[5]+tmp[7174]*kernel[6]+tmp[7175]*kernel[7]+tmp[7176]*kernel[8];
				ans[7076]<=tmp[6975]*kernel[0]+tmp[6976]*kernel[1]+tmp[6977]*kernel[2]+tmp[7075]*kernel[3]+tmp[7076]*kernel[4]+tmp[7077]*kernel[5]+tmp[7175]*kernel[6]+tmp[7176]*kernel[7]+tmp[7177]*kernel[8];
				ans[7077]<=tmp[6976]*kernel[0]+tmp[6977]*kernel[1]+tmp[6978]*kernel[2]+tmp[7076]*kernel[3]+tmp[7077]*kernel[4]+tmp[7078]*kernel[5]+tmp[7176]*kernel[6]+tmp[7177]*kernel[7]+tmp[7178]*kernel[8];
				ans[7078]<=tmp[6977]*kernel[0]+tmp[6978]*kernel[1]+tmp[6979]*kernel[2]+tmp[7077]*kernel[3]+tmp[7078]*kernel[4]+tmp[7079]*kernel[5]+tmp[7177]*kernel[6]+tmp[7178]*kernel[7]+tmp[7179]*kernel[8];
				ans[7079]<=tmp[6978]*kernel[0]+tmp[6979]*kernel[1]+tmp[6980]*kernel[2]+tmp[7078]*kernel[3]+tmp[7079]*kernel[4]+tmp[7080]*kernel[5]+tmp[7178]*kernel[6]+tmp[7179]*kernel[7]+tmp[7180]*kernel[8];
				ans[7080]<=tmp[6979]*kernel[0]+tmp[6980]*kernel[1]+tmp[6981]*kernel[2]+tmp[7079]*kernel[3]+tmp[7080]*kernel[4]+tmp[7081]*kernel[5]+tmp[7179]*kernel[6]+tmp[7180]*kernel[7]+tmp[7181]*kernel[8];
				ans[7081]<=tmp[6980]*kernel[0]+tmp[6981]*kernel[1]+tmp[6982]*kernel[2]+tmp[7080]*kernel[3]+tmp[7081]*kernel[4]+tmp[7082]*kernel[5]+tmp[7180]*kernel[6]+tmp[7181]*kernel[7]+tmp[7182]*kernel[8];
				ans[7082]<=tmp[6981]*kernel[0]+tmp[6982]*kernel[1]+tmp[6983]*kernel[2]+tmp[7081]*kernel[3]+tmp[7082]*kernel[4]+tmp[7083]*kernel[5]+tmp[7181]*kernel[6]+tmp[7182]*kernel[7]+tmp[7183]*kernel[8];
				ans[7083]<=tmp[6982]*kernel[0]+tmp[6983]*kernel[1]+tmp[6984]*kernel[2]+tmp[7082]*kernel[3]+tmp[7083]*kernel[4]+tmp[7084]*kernel[5]+tmp[7182]*kernel[6]+tmp[7183]*kernel[7]+tmp[7184]*kernel[8];
				ans[7084]<=tmp[6983]*kernel[0]+tmp[6984]*kernel[1]+tmp[6985]*kernel[2]+tmp[7083]*kernel[3]+tmp[7084]*kernel[4]+tmp[7085]*kernel[5]+tmp[7183]*kernel[6]+tmp[7184]*kernel[7]+tmp[7185]*kernel[8];
				ans[7085]<=tmp[6984]*kernel[0]+tmp[6985]*kernel[1]+tmp[6986]*kernel[2]+tmp[7084]*kernel[3]+tmp[7085]*kernel[4]+tmp[7086]*kernel[5]+tmp[7184]*kernel[6]+tmp[7185]*kernel[7]+tmp[7186]*kernel[8];
				ans[7086]<=tmp[6985]*kernel[0]+tmp[6986]*kernel[1]+tmp[6987]*kernel[2]+tmp[7085]*kernel[3]+tmp[7086]*kernel[4]+tmp[7087]*kernel[5]+tmp[7185]*kernel[6]+tmp[7186]*kernel[7]+tmp[7187]*kernel[8];
				ans[7087]<=tmp[6986]*kernel[0]+tmp[6987]*kernel[1]+tmp[6988]*kernel[2]+tmp[7086]*kernel[3]+tmp[7087]*kernel[4]+tmp[7088]*kernel[5]+tmp[7186]*kernel[6]+tmp[7187]*kernel[7]+tmp[7188]*kernel[8];
				ans[7088]<=tmp[6987]*kernel[0]+tmp[6988]*kernel[1]+tmp[6989]*kernel[2]+tmp[7087]*kernel[3]+tmp[7088]*kernel[4]+tmp[7089]*kernel[5]+tmp[7187]*kernel[6]+tmp[7188]*kernel[7]+tmp[7189]*kernel[8];
				ans[7089]<=tmp[6988]*kernel[0]+tmp[6989]*kernel[1]+tmp[6990]*kernel[2]+tmp[7088]*kernel[3]+tmp[7089]*kernel[4]+tmp[7090]*kernel[5]+tmp[7188]*kernel[6]+tmp[7189]*kernel[7]+tmp[7190]*kernel[8];
				ans[7090]<=tmp[6989]*kernel[0]+tmp[6990]*kernel[1]+tmp[6991]*kernel[2]+tmp[7089]*kernel[3]+tmp[7090]*kernel[4]+tmp[7091]*kernel[5]+tmp[7189]*kernel[6]+tmp[7190]*kernel[7]+tmp[7191]*kernel[8];
				ans[7091]<=tmp[6990]*kernel[0]+tmp[6991]*kernel[1]+tmp[6992]*kernel[2]+tmp[7090]*kernel[3]+tmp[7091]*kernel[4]+tmp[7092]*kernel[5]+tmp[7190]*kernel[6]+tmp[7191]*kernel[7]+tmp[7192]*kernel[8];
				ans[7092]<=tmp[6991]*kernel[0]+tmp[6992]*kernel[1]+tmp[6993]*kernel[2]+tmp[7091]*kernel[3]+tmp[7092]*kernel[4]+tmp[7093]*kernel[5]+tmp[7191]*kernel[6]+tmp[7192]*kernel[7]+tmp[7193]*kernel[8];
				ans[7093]<=tmp[6992]*kernel[0]+tmp[6993]*kernel[1]+tmp[6994]*kernel[2]+tmp[7092]*kernel[3]+tmp[7093]*kernel[4]+tmp[7094]*kernel[5]+tmp[7192]*kernel[6]+tmp[7193]*kernel[7]+tmp[7194]*kernel[8];
				ans[7094]<=tmp[6993]*kernel[0]+tmp[6994]*kernel[1]+tmp[6995]*kernel[2]+tmp[7093]*kernel[3]+tmp[7094]*kernel[4]+tmp[7095]*kernel[5]+tmp[7193]*kernel[6]+tmp[7194]*kernel[7]+tmp[7195]*kernel[8];
				ans[7095]<=tmp[6994]*kernel[0]+tmp[6995]*kernel[1]+tmp[6996]*kernel[2]+tmp[7094]*kernel[3]+tmp[7095]*kernel[4]+tmp[7096]*kernel[5]+tmp[7194]*kernel[6]+tmp[7195]*kernel[7]+tmp[7196]*kernel[8];
				ans[7096]<=tmp[6995]*kernel[0]+tmp[6996]*kernel[1]+tmp[6997]*kernel[2]+tmp[7095]*kernel[3]+tmp[7096]*kernel[4]+tmp[7097]*kernel[5]+tmp[7195]*kernel[6]+tmp[7196]*kernel[7]+tmp[7197]*kernel[8];
				ans[7097]<=tmp[6996]*kernel[0]+tmp[6997]*kernel[1]+tmp[6998]*kernel[2]+tmp[7096]*kernel[3]+tmp[7097]*kernel[4]+tmp[7098]*kernel[5]+tmp[7196]*kernel[6]+tmp[7197]*kernel[7]+tmp[7198]*kernel[8];
				ans[7098]<=tmp[6997]*kernel[0]+tmp[6998]*kernel[1]+tmp[6999]*kernel[2]+tmp[7097]*kernel[3]+tmp[7098]*kernel[4]+tmp[7099]*kernel[5]+tmp[7197]*kernel[6]+tmp[7198]*kernel[7]+tmp[7199]*kernel[8];
				ans[7099]<=tmp[6998]*kernel[0]+tmp[6999]*kernel[1]+tmp[7098]*kernel[3]+tmp[7099]*kernel[4]+tmp[7198]*kernel[6]+tmp[7199]*kernel[7];
				ans[7100]<=tmp[7000]*kernel[1]+tmp[7001]*kernel[2]+tmp[7100]*kernel[4]+tmp[7101]*kernel[5]+tmp[7200]*kernel[7]+tmp[7201]*kernel[8];
				ans[7101]<=tmp[7000]*kernel[0]+tmp[7001]*kernel[1]+tmp[7002]*kernel[2]+tmp[7100]*kernel[3]+tmp[7101]*kernel[4]+tmp[7102]*kernel[5]+tmp[7200]*kernel[6]+tmp[7201]*kernel[7]+tmp[7202]*kernel[8];
				ans[7102]<=tmp[7001]*kernel[0]+tmp[7002]*kernel[1]+tmp[7003]*kernel[2]+tmp[7101]*kernel[3]+tmp[7102]*kernel[4]+tmp[7103]*kernel[5]+tmp[7201]*kernel[6]+tmp[7202]*kernel[7]+tmp[7203]*kernel[8];
				ans[7103]<=tmp[7002]*kernel[0]+tmp[7003]*kernel[1]+tmp[7004]*kernel[2]+tmp[7102]*kernel[3]+tmp[7103]*kernel[4]+tmp[7104]*kernel[5]+tmp[7202]*kernel[6]+tmp[7203]*kernel[7]+tmp[7204]*kernel[8];
				ans[7104]<=tmp[7003]*kernel[0]+tmp[7004]*kernel[1]+tmp[7005]*kernel[2]+tmp[7103]*kernel[3]+tmp[7104]*kernel[4]+tmp[7105]*kernel[5]+tmp[7203]*kernel[6]+tmp[7204]*kernel[7]+tmp[7205]*kernel[8];
				ans[7105]<=tmp[7004]*kernel[0]+tmp[7005]*kernel[1]+tmp[7006]*kernel[2]+tmp[7104]*kernel[3]+tmp[7105]*kernel[4]+tmp[7106]*kernel[5]+tmp[7204]*kernel[6]+tmp[7205]*kernel[7]+tmp[7206]*kernel[8];
				ans[7106]<=tmp[7005]*kernel[0]+tmp[7006]*kernel[1]+tmp[7007]*kernel[2]+tmp[7105]*kernel[3]+tmp[7106]*kernel[4]+tmp[7107]*kernel[5]+tmp[7205]*kernel[6]+tmp[7206]*kernel[7]+tmp[7207]*kernel[8];
				ans[7107]<=tmp[7006]*kernel[0]+tmp[7007]*kernel[1]+tmp[7008]*kernel[2]+tmp[7106]*kernel[3]+tmp[7107]*kernel[4]+tmp[7108]*kernel[5]+tmp[7206]*kernel[6]+tmp[7207]*kernel[7]+tmp[7208]*kernel[8];
				ans[7108]<=tmp[7007]*kernel[0]+tmp[7008]*kernel[1]+tmp[7009]*kernel[2]+tmp[7107]*kernel[3]+tmp[7108]*kernel[4]+tmp[7109]*kernel[5]+tmp[7207]*kernel[6]+tmp[7208]*kernel[7]+tmp[7209]*kernel[8];
				ans[7109]<=tmp[7008]*kernel[0]+tmp[7009]*kernel[1]+tmp[7010]*kernel[2]+tmp[7108]*kernel[3]+tmp[7109]*kernel[4]+tmp[7110]*kernel[5]+tmp[7208]*kernel[6]+tmp[7209]*kernel[7]+tmp[7210]*kernel[8];
				ans[7110]<=tmp[7009]*kernel[0]+tmp[7010]*kernel[1]+tmp[7011]*kernel[2]+tmp[7109]*kernel[3]+tmp[7110]*kernel[4]+tmp[7111]*kernel[5]+tmp[7209]*kernel[6]+tmp[7210]*kernel[7]+tmp[7211]*kernel[8];
				ans[7111]<=tmp[7010]*kernel[0]+tmp[7011]*kernel[1]+tmp[7012]*kernel[2]+tmp[7110]*kernel[3]+tmp[7111]*kernel[4]+tmp[7112]*kernel[5]+tmp[7210]*kernel[6]+tmp[7211]*kernel[7]+tmp[7212]*kernel[8];
				ans[7112]<=tmp[7011]*kernel[0]+tmp[7012]*kernel[1]+tmp[7013]*kernel[2]+tmp[7111]*kernel[3]+tmp[7112]*kernel[4]+tmp[7113]*kernel[5]+tmp[7211]*kernel[6]+tmp[7212]*kernel[7]+tmp[7213]*kernel[8];
				ans[7113]<=tmp[7012]*kernel[0]+tmp[7013]*kernel[1]+tmp[7014]*kernel[2]+tmp[7112]*kernel[3]+tmp[7113]*kernel[4]+tmp[7114]*kernel[5]+tmp[7212]*kernel[6]+tmp[7213]*kernel[7]+tmp[7214]*kernel[8];
				ans[7114]<=tmp[7013]*kernel[0]+tmp[7014]*kernel[1]+tmp[7015]*kernel[2]+tmp[7113]*kernel[3]+tmp[7114]*kernel[4]+tmp[7115]*kernel[5]+tmp[7213]*kernel[6]+tmp[7214]*kernel[7]+tmp[7215]*kernel[8];
				ans[7115]<=tmp[7014]*kernel[0]+tmp[7015]*kernel[1]+tmp[7016]*kernel[2]+tmp[7114]*kernel[3]+tmp[7115]*kernel[4]+tmp[7116]*kernel[5]+tmp[7214]*kernel[6]+tmp[7215]*kernel[7]+tmp[7216]*kernel[8];
				ans[7116]<=tmp[7015]*kernel[0]+tmp[7016]*kernel[1]+tmp[7017]*kernel[2]+tmp[7115]*kernel[3]+tmp[7116]*kernel[4]+tmp[7117]*kernel[5]+tmp[7215]*kernel[6]+tmp[7216]*kernel[7]+tmp[7217]*kernel[8];
				ans[7117]<=tmp[7016]*kernel[0]+tmp[7017]*kernel[1]+tmp[7018]*kernel[2]+tmp[7116]*kernel[3]+tmp[7117]*kernel[4]+tmp[7118]*kernel[5]+tmp[7216]*kernel[6]+tmp[7217]*kernel[7]+tmp[7218]*kernel[8];
				ans[7118]<=tmp[7017]*kernel[0]+tmp[7018]*kernel[1]+tmp[7019]*kernel[2]+tmp[7117]*kernel[3]+tmp[7118]*kernel[4]+tmp[7119]*kernel[5]+tmp[7217]*kernel[6]+tmp[7218]*kernel[7]+tmp[7219]*kernel[8];
				ans[7119]<=tmp[7018]*kernel[0]+tmp[7019]*kernel[1]+tmp[7020]*kernel[2]+tmp[7118]*kernel[3]+tmp[7119]*kernel[4]+tmp[7120]*kernel[5]+tmp[7218]*kernel[6]+tmp[7219]*kernel[7]+tmp[7220]*kernel[8];
				ans[7120]<=tmp[7019]*kernel[0]+tmp[7020]*kernel[1]+tmp[7021]*kernel[2]+tmp[7119]*kernel[3]+tmp[7120]*kernel[4]+tmp[7121]*kernel[5]+tmp[7219]*kernel[6]+tmp[7220]*kernel[7]+tmp[7221]*kernel[8];
				ans[7121]<=tmp[7020]*kernel[0]+tmp[7021]*kernel[1]+tmp[7022]*kernel[2]+tmp[7120]*kernel[3]+tmp[7121]*kernel[4]+tmp[7122]*kernel[5]+tmp[7220]*kernel[6]+tmp[7221]*kernel[7]+tmp[7222]*kernel[8];
				ans[7122]<=tmp[7021]*kernel[0]+tmp[7022]*kernel[1]+tmp[7023]*kernel[2]+tmp[7121]*kernel[3]+tmp[7122]*kernel[4]+tmp[7123]*kernel[5]+tmp[7221]*kernel[6]+tmp[7222]*kernel[7]+tmp[7223]*kernel[8];
				ans[7123]<=tmp[7022]*kernel[0]+tmp[7023]*kernel[1]+tmp[7024]*kernel[2]+tmp[7122]*kernel[3]+tmp[7123]*kernel[4]+tmp[7124]*kernel[5]+tmp[7222]*kernel[6]+tmp[7223]*kernel[7]+tmp[7224]*kernel[8];
				ans[7124]<=tmp[7023]*kernel[0]+tmp[7024]*kernel[1]+tmp[7025]*kernel[2]+tmp[7123]*kernel[3]+tmp[7124]*kernel[4]+tmp[7125]*kernel[5]+tmp[7223]*kernel[6]+tmp[7224]*kernel[7]+tmp[7225]*kernel[8];
				ans[7125]<=tmp[7024]*kernel[0]+tmp[7025]*kernel[1]+tmp[7026]*kernel[2]+tmp[7124]*kernel[3]+tmp[7125]*kernel[4]+tmp[7126]*kernel[5]+tmp[7224]*kernel[6]+tmp[7225]*kernel[7]+tmp[7226]*kernel[8];
				ans[7126]<=tmp[7025]*kernel[0]+tmp[7026]*kernel[1]+tmp[7027]*kernel[2]+tmp[7125]*kernel[3]+tmp[7126]*kernel[4]+tmp[7127]*kernel[5]+tmp[7225]*kernel[6]+tmp[7226]*kernel[7]+tmp[7227]*kernel[8];
				ans[7127]<=tmp[7026]*kernel[0]+tmp[7027]*kernel[1]+tmp[7028]*kernel[2]+tmp[7126]*kernel[3]+tmp[7127]*kernel[4]+tmp[7128]*kernel[5]+tmp[7226]*kernel[6]+tmp[7227]*kernel[7]+tmp[7228]*kernel[8];
				ans[7128]<=tmp[7027]*kernel[0]+tmp[7028]*kernel[1]+tmp[7029]*kernel[2]+tmp[7127]*kernel[3]+tmp[7128]*kernel[4]+tmp[7129]*kernel[5]+tmp[7227]*kernel[6]+tmp[7228]*kernel[7]+tmp[7229]*kernel[8];
				ans[7129]<=tmp[7028]*kernel[0]+tmp[7029]*kernel[1]+tmp[7030]*kernel[2]+tmp[7128]*kernel[3]+tmp[7129]*kernel[4]+tmp[7130]*kernel[5]+tmp[7228]*kernel[6]+tmp[7229]*kernel[7]+tmp[7230]*kernel[8];
				ans[7130]<=tmp[7029]*kernel[0]+tmp[7030]*kernel[1]+tmp[7031]*kernel[2]+tmp[7129]*kernel[3]+tmp[7130]*kernel[4]+tmp[7131]*kernel[5]+tmp[7229]*kernel[6]+tmp[7230]*kernel[7]+tmp[7231]*kernel[8];
				ans[7131]<=tmp[7030]*kernel[0]+tmp[7031]*kernel[1]+tmp[7032]*kernel[2]+tmp[7130]*kernel[3]+tmp[7131]*kernel[4]+tmp[7132]*kernel[5]+tmp[7230]*kernel[6]+tmp[7231]*kernel[7]+tmp[7232]*kernel[8];
				ans[7132]<=tmp[7031]*kernel[0]+tmp[7032]*kernel[1]+tmp[7033]*kernel[2]+tmp[7131]*kernel[3]+tmp[7132]*kernel[4]+tmp[7133]*kernel[5]+tmp[7231]*kernel[6]+tmp[7232]*kernel[7]+tmp[7233]*kernel[8];
				ans[7133]<=tmp[7032]*kernel[0]+tmp[7033]*kernel[1]+tmp[7034]*kernel[2]+tmp[7132]*kernel[3]+tmp[7133]*kernel[4]+tmp[7134]*kernel[5]+tmp[7232]*kernel[6]+tmp[7233]*kernel[7]+tmp[7234]*kernel[8];
				ans[7134]<=tmp[7033]*kernel[0]+tmp[7034]*kernel[1]+tmp[7035]*kernel[2]+tmp[7133]*kernel[3]+tmp[7134]*kernel[4]+tmp[7135]*kernel[5]+tmp[7233]*kernel[6]+tmp[7234]*kernel[7]+tmp[7235]*kernel[8];
				ans[7135]<=tmp[7034]*kernel[0]+tmp[7035]*kernel[1]+tmp[7036]*kernel[2]+tmp[7134]*kernel[3]+tmp[7135]*kernel[4]+tmp[7136]*kernel[5]+tmp[7234]*kernel[6]+tmp[7235]*kernel[7]+tmp[7236]*kernel[8];
				ans[7136]<=tmp[7035]*kernel[0]+tmp[7036]*kernel[1]+tmp[7037]*kernel[2]+tmp[7135]*kernel[3]+tmp[7136]*kernel[4]+tmp[7137]*kernel[5]+tmp[7235]*kernel[6]+tmp[7236]*kernel[7]+tmp[7237]*kernel[8];
				ans[7137]<=tmp[7036]*kernel[0]+tmp[7037]*kernel[1]+tmp[7038]*kernel[2]+tmp[7136]*kernel[3]+tmp[7137]*kernel[4]+tmp[7138]*kernel[5]+tmp[7236]*kernel[6]+tmp[7237]*kernel[7]+tmp[7238]*kernel[8];
				ans[7138]<=tmp[7037]*kernel[0]+tmp[7038]*kernel[1]+tmp[7039]*kernel[2]+tmp[7137]*kernel[3]+tmp[7138]*kernel[4]+tmp[7139]*kernel[5]+tmp[7237]*kernel[6]+tmp[7238]*kernel[7]+tmp[7239]*kernel[8];
				ans[7139]<=tmp[7038]*kernel[0]+tmp[7039]*kernel[1]+tmp[7040]*kernel[2]+tmp[7138]*kernel[3]+tmp[7139]*kernel[4]+tmp[7140]*kernel[5]+tmp[7238]*kernel[6]+tmp[7239]*kernel[7]+tmp[7240]*kernel[8];
				ans[7140]<=tmp[7039]*kernel[0]+tmp[7040]*kernel[1]+tmp[7041]*kernel[2]+tmp[7139]*kernel[3]+tmp[7140]*kernel[4]+tmp[7141]*kernel[5]+tmp[7239]*kernel[6]+tmp[7240]*kernel[7]+tmp[7241]*kernel[8];
				ans[7141]<=tmp[7040]*kernel[0]+tmp[7041]*kernel[1]+tmp[7042]*kernel[2]+tmp[7140]*kernel[3]+tmp[7141]*kernel[4]+tmp[7142]*kernel[5]+tmp[7240]*kernel[6]+tmp[7241]*kernel[7]+tmp[7242]*kernel[8];
				ans[7142]<=tmp[7041]*kernel[0]+tmp[7042]*kernel[1]+tmp[7043]*kernel[2]+tmp[7141]*kernel[3]+tmp[7142]*kernel[4]+tmp[7143]*kernel[5]+tmp[7241]*kernel[6]+tmp[7242]*kernel[7]+tmp[7243]*kernel[8];
				ans[7143]<=tmp[7042]*kernel[0]+tmp[7043]*kernel[1]+tmp[7044]*kernel[2]+tmp[7142]*kernel[3]+tmp[7143]*kernel[4]+tmp[7144]*kernel[5]+tmp[7242]*kernel[6]+tmp[7243]*kernel[7]+tmp[7244]*kernel[8];
				ans[7144]<=tmp[7043]*kernel[0]+tmp[7044]*kernel[1]+tmp[7045]*kernel[2]+tmp[7143]*kernel[3]+tmp[7144]*kernel[4]+tmp[7145]*kernel[5]+tmp[7243]*kernel[6]+tmp[7244]*kernel[7]+tmp[7245]*kernel[8];
				ans[7145]<=tmp[7044]*kernel[0]+tmp[7045]*kernel[1]+tmp[7046]*kernel[2]+tmp[7144]*kernel[3]+tmp[7145]*kernel[4]+tmp[7146]*kernel[5]+tmp[7244]*kernel[6]+tmp[7245]*kernel[7]+tmp[7246]*kernel[8];
				ans[7146]<=tmp[7045]*kernel[0]+tmp[7046]*kernel[1]+tmp[7047]*kernel[2]+tmp[7145]*kernel[3]+tmp[7146]*kernel[4]+tmp[7147]*kernel[5]+tmp[7245]*kernel[6]+tmp[7246]*kernel[7]+tmp[7247]*kernel[8];
				ans[7147]<=tmp[7046]*kernel[0]+tmp[7047]*kernel[1]+tmp[7048]*kernel[2]+tmp[7146]*kernel[3]+tmp[7147]*kernel[4]+tmp[7148]*kernel[5]+tmp[7246]*kernel[6]+tmp[7247]*kernel[7]+tmp[7248]*kernel[8];
				ans[7148]<=tmp[7047]*kernel[0]+tmp[7048]*kernel[1]+tmp[7049]*kernel[2]+tmp[7147]*kernel[3]+tmp[7148]*kernel[4]+tmp[7149]*kernel[5]+tmp[7247]*kernel[6]+tmp[7248]*kernel[7]+tmp[7249]*kernel[8];
				ans[7149]<=tmp[7048]*kernel[0]+tmp[7049]*kernel[1]+tmp[7050]*kernel[2]+tmp[7148]*kernel[3]+tmp[7149]*kernel[4]+tmp[7150]*kernel[5]+tmp[7248]*kernel[6]+tmp[7249]*kernel[7]+tmp[7250]*kernel[8];
				ans[7150]<=tmp[7049]*kernel[0]+tmp[7050]*kernel[1]+tmp[7051]*kernel[2]+tmp[7149]*kernel[3]+tmp[7150]*kernel[4]+tmp[7151]*kernel[5]+tmp[7249]*kernel[6]+tmp[7250]*kernel[7]+tmp[7251]*kernel[8];
				ans[7151]<=tmp[7050]*kernel[0]+tmp[7051]*kernel[1]+tmp[7052]*kernel[2]+tmp[7150]*kernel[3]+tmp[7151]*kernel[4]+tmp[7152]*kernel[5]+tmp[7250]*kernel[6]+tmp[7251]*kernel[7]+tmp[7252]*kernel[8];
				ans[7152]<=tmp[7051]*kernel[0]+tmp[7052]*kernel[1]+tmp[7053]*kernel[2]+tmp[7151]*kernel[3]+tmp[7152]*kernel[4]+tmp[7153]*kernel[5]+tmp[7251]*kernel[6]+tmp[7252]*kernel[7]+tmp[7253]*kernel[8];
				ans[7153]<=tmp[7052]*kernel[0]+tmp[7053]*kernel[1]+tmp[7054]*kernel[2]+tmp[7152]*kernel[3]+tmp[7153]*kernel[4]+tmp[7154]*kernel[5]+tmp[7252]*kernel[6]+tmp[7253]*kernel[7]+tmp[7254]*kernel[8];
				ans[7154]<=tmp[7053]*kernel[0]+tmp[7054]*kernel[1]+tmp[7055]*kernel[2]+tmp[7153]*kernel[3]+tmp[7154]*kernel[4]+tmp[7155]*kernel[5]+tmp[7253]*kernel[6]+tmp[7254]*kernel[7]+tmp[7255]*kernel[8];
				ans[7155]<=tmp[7054]*kernel[0]+tmp[7055]*kernel[1]+tmp[7056]*kernel[2]+tmp[7154]*kernel[3]+tmp[7155]*kernel[4]+tmp[7156]*kernel[5]+tmp[7254]*kernel[6]+tmp[7255]*kernel[7]+tmp[7256]*kernel[8];
				ans[7156]<=tmp[7055]*kernel[0]+tmp[7056]*kernel[1]+tmp[7057]*kernel[2]+tmp[7155]*kernel[3]+tmp[7156]*kernel[4]+tmp[7157]*kernel[5]+tmp[7255]*kernel[6]+tmp[7256]*kernel[7]+tmp[7257]*kernel[8];
				ans[7157]<=tmp[7056]*kernel[0]+tmp[7057]*kernel[1]+tmp[7058]*kernel[2]+tmp[7156]*kernel[3]+tmp[7157]*kernel[4]+tmp[7158]*kernel[5]+tmp[7256]*kernel[6]+tmp[7257]*kernel[7]+tmp[7258]*kernel[8];
				ans[7158]<=tmp[7057]*kernel[0]+tmp[7058]*kernel[1]+tmp[7059]*kernel[2]+tmp[7157]*kernel[3]+tmp[7158]*kernel[4]+tmp[7159]*kernel[5]+tmp[7257]*kernel[6]+tmp[7258]*kernel[7]+tmp[7259]*kernel[8];
				ans[7159]<=tmp[7058]*kernel[0]+tmp[7059]*kernel[1]+tmp[7060]*kernel[2]+tmp[7158]*kernel[3]+tmp[7159]*kernel[4]+tmp[7160]*kernel[5]+tmp[7258]*kernel[6]+tmp[7259]*kernel[7]+tmp[7260]*kernel[8];
				ans[7160]<=tmp[7059]*kernel[0]+tmp[7060]*kernel[1]+tmp[7061]*kernel[2]+tmp[7159]*kernel[3]+tmp[7160]*kernel[4]+tmp[7161]*kernel[5]+tmp[7259]*kernel[6]+tmp[7260]*kernel[7]+tmp[7261]*kernel[8];
				ans[7161]<=tmp[7060]*kernel[0]+tmp[7061]*kernel[1]+tmp[7062]*kernel[2]+tmp[7160]*kernel[3]+tmp[7161]*kernel[4]+tmp[7162]*kernel[5]+tmp[7260]*kernel[6]+tmp[7261]*kernel[7]+tmp[7262]*kernel[8];
				ans[7162]<=tmp[7061]*kernel[0]+tmp[7062]*kernel[1]+tmp[7063]*kernel[2]+tmp[7161]*kernel[3]+tmp[7162]*kernel[4]+tmp[7163]*kernel[5]+tmp[7261]*kernel[6]+tmp[7262]*kernel[7]+tmp[7263]*kernel[8];
				ans[7163]<=tmp[7062]*kernel[0]+tmp[7063]*kernel[1]+tmp[7064]*kernel[2]+tmp[7162]*kernel[3]+tmp[7163]*kernel[4]+tmp[7164]*kernel[5]+tmp[7262]*kernel[6]+tmp[7263]*kernel[7]+tmp[7264]*kernel[8];
				ans[7164]<=tmp[7063]*kernel[0]+tmp[7064]*kernel[1]+tmp[7065]*kernel[2]+tmp[7163]*kernel[3]+tmp[7164]*kernel[4]+tmp[7165]*kernel[5]+tmp[7263]*kernel[6]+tmp[7264]*kernel[7]+tmp[7265]*kernel[8];
				ans[7165]<=tmp[7064]*kernel[0]+tmp[7065]*kernel[1]+tmp[7066]*kernel[2]+tmp[7164]*kernel[3]+tmp[7165]*kernel[4]+tmp[7166]*kernel[5]+tmp[7264]*kernel[6]+tmp[7265]*kernel[7]+tmp[7266]*kernel[8];
				ans[7166]<=tmp[7065]*kernel[0]+tmp[7066]*kernel[1]+tmp[7067]*kernel[2]+tmp[7165]*kernel[3]+tmp[7166]*kernel[4]+tmp[7167]*kernel[5]+tmp[7265]*kernel[6]+tmp[7266]*kernel[7]+tmp[7267]*kernel[8];
				ans[7167]<=tmp[7066]*kernel[0]+tmp[7067]*kernel[1]+tmp[7068]*kernel[2]+tmp[7166]*kernel[3]+tmp[7167]*kernel[4]+tmp[7168]*kernel[5]+tmp[7266]*kernel[6]+tmp[7267]*kernel[7]+tmp[7268]*kernel[8];
				ans[7168]<=tmp[7067]*kernel[0]+tmp[7068]*kernel[1]+tmp[7069]*kernel[2]+tmp[7167]*kernel[3]+tmp[7168]*kernel[4]+tmp[7169]*kernel[5]+tmp[7267]*kernel[6]+tmp[7268]*kernel[7]+tmp[7269]*kernel[8];
				ans[7169]<=tmp[7068]*kernel[0]+tmp[7069]*kernel[1]+tmp[7070]*kernel[2]+tmp[7168]*kernel[3]+tmp[7169]*kernel[4]+tmp[7170]*kernel[5]+tmp[7268]*kernel[6]+tmp[7269]*kernel[7]+tmp[7270]*kernel[8];
				ans[7170]<=tmp[7069]*kernel[0]+tmp[7070]*kernel[1]+tmp[7071]*kernel[2]+tmp[7169]*kernel[3]+tmp[7170]*kernel[4]+tmp[7171]*kernel[5]+tmp[7269]*kernel[6]+tmp[7270]*kernel[7]+tmp[7271]*kernel[8];
				ans[7171]<=tmp[7070]*kernel[0]+tmp[7071]*kernel[1]+tmp[7072]*kernel[2]+tmp[7170]*kernel[3]+tmp[7171]*kernel[4]+tmp[7172]*kernel[5]+tmp[7270]*kernel[6]+tmp[7271]*kernel[7]+tmp[7272]*kernel[8];
				ans[7172]<=tmp[7071]*kernel[0]+tmp[7072]*kernel[1]+tmp[7073]*kernel[2]+tmp[7171]*kernel[3]+tmp[7172]*kernel[4]+tmp[7173]*kernel[5]+tmp[7271]*kernel[6]+tmp[7272]*kernel[7]+tmp[7273]*kernel[8];
				ans[7173]<=tmp[7072]*kernel[0]+tmp[7073]*kernel[1]+tmp[7074]*kernel[2]+tmp[7172]*kernel[3]+tmp[7173]*kernel[4]+tmp[7174]*kernel[5]+tmp[7272]*kernel[6]+tmp[7273]*kernel[7]+tmp[7274]*kernel[8];
				ans[7174]<=tmp[7073]*kernel[0]+tmp[7074]*kernel[1]+tmp[7075]*kernel[2]+tmp[7173]*kernel[3]+tmp[7174]*kernel[4]+tmp[7175]*kernel[5]+tmp[7273]*kernel[6]+tmp[7274]*kernel[7]+tmp[7275]*kernel[8];
				ans[7175]<=tmp[7074]*kernel[0]+tmp[7075]*kernel[1]+tmp[7076]*kernel[2]+tmp[7174]*kernel[3]+tmp[7175]*kernel[4]+tmp[7176]*kernel[5]+tmp[7274]*kernel[6]+tmp[7275]*kernel[7]+tmp[7276]*kernel[8];
				ans[7176]<=tmp[7075]*kernel[0]+tmp[7076]*kernel[1]+tmp[7077]*kernel[2]+tmp[7175]*kernel[3]+tmp[7176]*kernel[4]+tmp[7177]*kernel[5]+tmp[7275]*kernel[6]+tmp[7276]*kernel[7]+tmp[7277]*kernel[8];
				ans[7177]<=tmp[7076]*kernel[0]+tmp[7077]*kernel[1]+tmp[7078]*kernel[2]+tmp[7176]*kernel[3]+tmp[7177]*kernel[4]+tmp[7178]*kernel[5]+tmp[7276]*kernel[6]+tmp[7277]*kernel[7]+tmp[7278]*kernel[8];
				ans[7178]<=tmp[7077]*kernel[0]+tmp[7078]*kernel[1]+tmp[7079]*kernel[2]+tmp[7177]*kernel[3]+tmp[7178]*kernel[4]+tmp[7179]*kernel[5]+tmp[7277]*kernel[6]+tmp[7278]*kernel[7]+tmp[7279]*kernel[8];
				ans[7179]<=tmp[7078]*kernel[0]+tmp[7079]*kernel[1]+tmp[7080]*kernel[2]+tmp[7178]*kernel[3]+tmp[7179]*kernel[4]+tmp[7180]*kernel[5]+tmp[7278]*kernel[6]+tmp[7279]*kernel[7]+tmp[7280]*kernel[8];
				ans[7180]<=tmp[7079]*kernel[0]+tmp[7080]*kernel[1]+tmp[7081]*kernel[2]+tmp[7179]*kernel[3]+tmp[7180]*kernel[4]+tmp[7181]*kernel[5]+tmp[7279]*kernel[6]+tmp[7280]*kernel[7]+tmp[7281]*kernel[8];
				ans[7181]<=tmp[7080]*kernel[0]+tmp[7081]*kernel[1]+tmp[7082]*kernel[2]+tmp[7180]*kernel[3]+tmp[7181]*kernel[4]+tmp[7182]*kernel[5]+tmp[7280]*kernel[6]+tmp[7281]*kernel[7]+tmp[7282]*kernel[8];
				ans[7182]<=tmp[7081]*kernel[0]+tmp[7082]*kernel[1]+tmp[7083]*kernel[2]+tmp[7181]*kernel[3]+tmp[7182]*kernel[4]+tmp[7183]*kernel[5]+tmp[7281]*kernel[6]+tmp[7282]*kernel[7]+tmp[7283]*kernel[8];
				ans[7183]<=tmp[7082]*kernel[0]+tmp[7083]*kernel[1]+tmp[7084]*kernel[2]+tmp[7182]*kernel[3]+tmp[7183]*kernel[4]+tmp[7184]*kernel[5]+tmp[7282]*kernel[6]+tmp[7283]*kernel[7]+tmp[7284]*kernel[8];
				ans[7184]<=tmp[7083]*kernel[0]+tmp[7084]*kernel[1]+tmp[7085]*kernel[2]+tmp[7183]*kernel[3]+tmp[7184]*kernel[4]+tmp[7185]*kernel[5]+tmp[7283]*kernel[6]+tmp[7284]*kernel[7]+tmp[7285]*kernel[8];
				ans[7185]<=tmp[7084]*kernel[0]+tmp[7085]*kernel[1]+tmp[7086]*kernel[2]+tmp[7184]*kernel[3]+tmp[7185]*kernel[4]+tmp[7186]*kernel[5]+tmp[7284]*kernel[6]+tmp[7285]*kernel[7]+tmp[7286]*kernel[8];
				ans[7186]<=tmp[7085]*kernel[0]+tmp[7086]*kernel[1]+tmp[7087]*kernel[2]+tmp[7185]*kernel[3]+tmp[7186]*kernel[4]+tmp[7187]*kernel[5]+tmp[7285]*kernel[6]+tmp[7286]*kernel[7]+tmp[7287]*kernel[8];
				ans[7187]<=tmp[7086]*kernel[0]+tmp[7087]*kernel[1]+tmp[7088]*kernel[2]+tmp[7186]*kernel[3]+tmp[7187]*kernel[4]+tmp[7188]*kernel[5]+tmp[7286]*kernel[6]+tmp[7287]*kernel[7]+tmp[7288]*kernel[8];
				ans[7188]<=tmp[7087]*kernel[0]+tmp[7088]*kernel[1]+tmp[7089]*kernel[2]+tmp[7187]*kernel[3]+tmp[7188]*kernel[4]+tmp[7189]*kernel[5]+tmp[7287]*kernel[6]+tmp[7288]*kernel[7]+tmp[7289]*kernel[8];
				ans[7189]<=tmp[7088]*kernel[0]+tmp[7089]*kernel[1]+tmp[7090]*kernel[2]+tmp[7188]*kernel[3]+tmp[7189]*kernel[4]+tmp[7190]*kernel[5]+tmp[7288]*kernel[6]+tmp[7289]*kernel[7]+tmp[7290]*kernel[8];
				ans[7190]<=tmp[7089]*kernel[0]+tmp[7090]*kernel[1]+tmp[7091]*kernel[2]+tmp[7189]*kernel[3]+tmp[7190]*kernel[4]+tmp[7191]*kernel[5]+tmp[7289]*kernel[6]+tmp[7290]*kernel[7]+tmp[7291]*kernel[8];
				ans[7191]<=tmp[7090]*kernel[0]+tmp[7091]*kernel[1]+tmp[7092]*kernel[2]+tmp[7190]*kernel[3]+tmp[7191]*kernel[4]+tmp[7192]*kernel[5]+tmp[7290]*kernel[6]+tmp[7291]*kernel[7]+tmp[7292]*kernel[8];
				ans[7192]<=tmp[7091]*kernel[0]+tmp[7092]*kernel[1]+tmp[7093]*kernel[2]+tmp[7191]*kernel[3]+tmp[7192]*kernel[4]+tmp[7193]*kernel[5]+tmp[7291]*kernel[6]+tmp[7292]*kernel[7]+tmp[7293]*kernel[8];
				ans[7193]<=tmp[7092]*kernel[0]+tmp[7093]*kernel[1]+tmp[7094]*kernel[2]+tmp[7192]*kernel[3]+tmp[7193]*kernel[4]+tmp[7194]*kernel[5]+tmp[7292]*kernel[6]+tmp[7293]*kernel[7]+tmp[7294]*kernel[8];
				ans[7194]<=tmp[7093]*kernel[0]+tmp[7094]*kernel[1]+tmp[7095]*kernel[2]+tmp[7193]*kernel[3]+tmp[7194]*kernel[4]+tmp[7195]*kernel[5]+tmp[7293]*kernel[6]+tmp[7294]*kernel[7]+tmp[7295]*kernel[8];
				ans[7195]<=tmp[7094]*kernel[0]+tmp[7095]*kernel[1]+tmp[7096]*kernel[2]+tmp[7194]*kernel[3]+tmp[7195]*kernel[4]+tmp[7196]*kernel[5]+tmp[7294]*kernel[6]+tmp[7295]*kernel[7]+tmp[7296]*kernel[8];
				ans[7196]<=tmp[7095]*kernel[0]+tmp[7096]*kernel[1]+tmp[7097]*kernel[2]+tmp[7195]*kernel[3]+tmp[7196]*kernel[4]+tmp[7197]*kernel[5]+tmp[7295]*kernel[6]+tmp[7296]*kernel[7]+tmp[7297]*kernel[8];
				ans[7197]<=tmp[7096]*kernel[0]+tmp[7097]*kernel[1]+tmp[7098]*kernel[2]+tmp[7196]*kernel[3]+tmp[7197]*kernel[4]+tmp[7198]*kernel[5]+tmp[7296]*kernel[6]+tmp[7297]*kernel[7]+tmp[7298]*kernel[8];
				ans[7198]<=tmp[7097]*kernel[0]+tmp[7098]*kernel[1]+tmp[7099]*kernel[2]+tmp[7197]*kernel[3]+tmp[7198]*kernel[4]+tmp[7199]*kernel[5]+tmp[7297]*kernel[6]+tmp[7298]*kernel[7]+tmp[7299]*kernel[8];
				ans[7199]<=tmp[7098]*kernel[0]+tmp[7099]*kernel[1]+tmp[7198]*kernel[3]+tmp[7199]*kernel[4]+tmp[7298]*kernel[6]+tmp[7299]*kernel[7];
				ans[7200]<=tmp[7100]*kernel[1]+tmp[7101]*kernel[2]+tmp[7200]*kernel[4]+tmp[7201]*kernel[5]+tmp[7300]*kernel[7]+tmp[7301]*kernel[8];
				ans[7201]<=tmp[7100]*kernel[0]+tmp[7101]*kernel[1]+tmp[7102]*kernel[2]+tmp[7200]*kernel[3]+tmp[7201]*kernel[4]+tmp[7202]*kernel[5]+tmp[7300]*kernel[6]+tmp[7301]*kernel[7]+tmp[7302]*kernel[8];
				ans[7202]<=tmp[7101]*kernel[0]+tmp[7102]*kernel[1]+tmp[7103]*kernel[2]+tmp[7201]*kernel[3]+tmp[7202]*kernel[4]+tmp[7203]*kernel[5]+tmp[7301]*kernel[6]+tmp[7302]*kernel[7]+tmp[7303]*kernel[8];
				ans[7203]<=tmp[7102]*kernel[0]+tmp[7103]*kernel[1]+tmp[7104]*kernel[2]+tmp[7202]*kernel[3]+tmp[7203]*kernel[4]+tmp[7204]*kernel[5]+tmp[7302]*kernel[6]+tmp[7303]*kernel[7]+tmp[7304]*kernel[8];
				ans[7204]<=tmp[7103]*kernel[0]+tmp[7104]*kernel[1]+tmp[7105]*kernel[2]+tmp[7203]*kernel[3]+tmp[7204]*kernel[4]+tmp[7205]*kernel[5]+tmp[7303]*kernel[6]+tmp[7304]*kernel[7]+tmp[7305]*kernel[8];
				ans[7205]<=tmp[7104]*kernel[0]+tmp[7105]*kernel[1]+tmp[7106]*kernel[2]+tmp[7204]*kernel[3]+tmp[7205]*kernel[4]+tmp[7206]*kernel[5]+tmp[7304]*kernel[6]+tmp[7305]*kernel[7]+tmp[7306]*kernel[8];
				ans[7206]<=tmp[7105]*kernel[0]+tmp[7106]*kernel[1]+tmp[7107]*kernel[2]+tmp[7205]*kernel[3]+tmp[7206]*kernel[4]+tmp[7207]*kernel[5]+tmp[7305]*kernel[6]+tmp[7306]*kernel[7]+tmp[7307]*kernel[8];
				ans[7207]<=tmp[7106]*kernel[0]+tmp[7107]*kernel[1]+tmp[7108]*kernel[2]+tmp[7206]*kernel[3]+tmp[7207]*kernel[4]+tmp[7208]*kernel[5]+tmp[7306]*kernel[6]+tmp[7307]*kernel[7]+tmp[7308]*kernel[8];
				ans[7208]<=tmp[7107]*kernel[0]+tmp[7108]*kernel[1]+tmp[7109]*kernel[2]+tmp[7207]*kernel[3]+tmp[7208]*kernel[4]+tmp[7209]*kernel[5]+tmp[7307]*kernel[6]+tmp[7308]*kernel[7]+tmp[7309]*kernel[8];
				ans[7209]<=tmp[7108]*kernel[0]+tmp[7109]*kernel[1]+tmp[7110]*kernel[2]+tmp[7208]*kernel[3]+tmp[7209]*kernel[4]+tmp[7210]*kernel[5]+tmp[7308]*kernel[6]+tmp[7309]*kernel[7]+tmp[7310]*kernel[8];
				ans[7210]<=tmp[7109]*kernel[0]+tmp[7110]*kernel[1]+tmp[7111]*kernel[2]+tmp[7209]*kernel[3]+tmp[7210]*kernel[4]+tmp[7211]*kernel[5]+tmp[7309]*kernel[6]+tmp[7310]*kernel[7]+tmp[7311]*kernel[8];
				ans[7211]<=tmp[7110]*kernel[0]+tmp[7111]*kernel[1]+tmp[7112]*kernel[2]+tmp[7210]*kernel[3]+tmp[7211]*kernel[4]+tmp[7212]*kernel[5]+tmp[7310]*kernel[6]+tmp[7311]*kernel[7]+tmp[7312]*kernel[8];
				ans[7212]<=tmp[7111]*kernel[0]+tmp[7112]*kernel[1]+tmp[7113]*kernel[2]+tmp[7211]*kernel[3]+tmp[7212]*kernel[4]+tmp[7213]*kernel[5]+tmp[7311]*kernel[6]+tmp[7312]*kernel[7]+tmp[7313]*kernel[8];
				ans[7213]<=tmp[7112]*kernel[0]+tmp[7113]*kernel[1]+tmp[7114]*kernel[2]+tmp[7212]*kernel[3]+tmp[7213]*kernel[4]+tmp[7214]*kernel[5]+tmp[7312]*kernel[6]+tmp[7313]*kernel[7]+tmp[7314]*kernel[8];
				ans[7214]<=tmp[7113]*kernel[0]+tmp[7114]*kernel[1]+tmp[7115]*kernel[2]+tmp[7213]*kernel[3]+tmp[7214]*kernel[4]+tmp[7215]*kernel[5]+tmp[7313]*kernel[6]+tmp[7314]*kernel[7]+tmp[7315]*kernel[8];
				ans[7215]<=tmp[7114]*kernel[0]+tmp[7115]*kernel[1]+tmp[7116]*kernel[2]+tmp[7214]*kernel[3]+tmp[7215]*kernel[4]+tmp[7216]*kernel[5]+tmp[7314]*kernel[6]+tmp[7315]*kernel[7]+tmp[7316]*kernel[8];
				ans[7216]<=tmp[7115]*kernel[0]+tmp[7116]*kernel[1]+tmp[7117]*kernel[2]+tmp[7215]*kernel[3]+tmp[7216]*kernel[4]+tmp[7217]*kernel[5]+tmp[7315]*kernel[6]+tmp[7316]*kernel[7]+tmp[7317]*kernel[8];
				ans[7217]<=tmp[7116]*kernel[0]+tmp[7117]*kernel[1]+tmp[7118]*kernel[2]+tmp[7216]*kernel[3]+tmp[7217]*kernel[4]+tmp[7218]*kernel[5]+tmp[7316]*kernel[6]+tmp[7317]*kernel[7]+tmp[7318]*kernel[8];
				ans[7218]<=tmp[7117]*kernel[0]+tmp[7118]*kernel[1]+tmp[7119]*kernel[2]+tmp[7217]*kernel[3]+tmp[7218]*kernel[4]+tmp[7219]*kernel[5]+tmp[7317]*kernel[6]+tmp[7318]*kernel[7]+tmp[7319]*kernel[8];
				ans[7219]<=tmp[7118]*kernel[0]+tmp[7119]*kernel[1]+tmp[7120]*kernel[2]+tmp[7218]*kernel[3]+tmp[7219]*kernel[4]+tmp[7220]*kernel[5]+tmp[7318]*kernel[6]+tmp[7319]*kernel[7]+tmp[7320]*kernel[8];
				ans[7220]<=tmp[7119]*kernel[0]+tmp[7120]*kernel[1]+tmp[7121]*kernel[2]+tmp[7219]*kernel[3]+tmp[7220]*kernel[4]+tmp[7221]*kernel[5]+tmp[7319]*kernel[6]+tmp[7320]*kernel[7]+tmp[7321]*kernel[8];
				ans[7221]<=tmp[7120]*kernel[0]+tmp[7121]*kernel[1]+tmp[7122]*kernel[2]+tmp[7220]*kernel[3]+tmp[7221]*kernel[4]+tmp[7222]*kernel[5]+tmp[7320]*kernel[6]+tmp[7321]*kernel[7]+tmp[7322]*kernel[8];
				ans[7222]<=tmp[7121]*kernel[0]+tmp[7122]*kernel[1]+tmp[7123]*kernel[2]+tmp[7221]*kernel[3]+tmp[7222]*kernel[4]+tmp[7223]*kernel[5]+tmp[7321]*kernel[6]+tmp[7322]*kernel[7]+tmp[7323]*kernel[8];
				ans[7223]<=tmp[7122]*kernel[0]+tmp[7123]*kernel[1]+tmp[7124]*kernel[2]+tmp[7222]*kernel[3]+tmp[7223]*kernel[4]+tmp[7224]*kernel[5]+tmp[7322]*kernel[6]+tmp[7323]*kernel[7]+tmp[7324]*kernel[8];
				ans[7224]<=tmp[7123]*kernel[0]+tmp[7124]*kernel[1]+tmp[7125]*kernel[2]+tmp[7223]*kernel[3]+tmp[7224]*kernel[4]+tmp[7225]*kernel[5]+tmp[7323]*kernel[6]+tmp[7324]*kernel[7]+tmp[7325]*kernel[8];
				ans[7225]<=tmp[7124]*kernel[0]+tmp[7125]*kernel[1]+tmp[7126]*kernel[2]+tmp[7224]*kernel[3]+tmp[7225]*kernel[4]+tmp[7226]*kernel[5]+tmp[7324]*kernel[6]+tmp[7325]*kernel[7]+tmp[7326]*kernel[8];
				ans[7226]<=tmp[7125]*kernel[0]+tmp[7126]*kernel[1]+tmp[7127]*kernel[2]+tmp[7225]*kernel[3]+tmp[7226]*kernel[4]+tmp[7227]*kernel[5]+tmp[7325]*kernel[6]+tmp[7326]*kernel[7]+tmp[7327]*kernel[8];
				ans[7227]<=tmp[7126]*kernel[0]+tmp[7127]*kernel[1]+tmp[7128]*kernel[2]+tmp[7226]*kernel[3]+tmp[7227]*kernel[4]+tmp[7228]*kernel[5]+tmp[7326]*kernel[6]+tmp[7327]*kernel[7]+tmp[7328]*kernel[8];
				ans[7228]<=tmp[7127]*kernel[0]+tmp[7128]*kernel[1]+tmp[7129]*kernel[2]+tmp[7227]*kernel[3]+tmp[7228]*kernel[4]+tmp[7229]*kernel[5]+tmp[7327]*kernel[6]+tmp[7328]*kernel[7]+tmp[7329]*kernel[8];
				ans[7229]<=tmp[7128]*kernel[0]+tmp[7129]*kernel[1]+tmp[7130]*kernel[2]+tmp[7228]*kernel[3]+tmp[7229]*kernel[4]+tmp[7230]*kernel[5]+tmp[7328]*kernel[6]+tmp[7329]*kernel[7]+tmp[7330]*kernel[8];
				ans[7230]<=tmp[7129]*kernel[0]+tmp[7130]*kernel[1]+tmp[7131]*kernel[2]+tmp[7229]*kernel[3]+tmp[7230]*kernel[4]+tmp[7231]*kernel[5]+tmp[7329]*kernel[6]+tmp[7330]*kernel[7]+tmp[7331]*kernel[8];
				ans[7231]<=tmp[7130]*kernel[0]+tmp[7131]*kernel[1]+tmp[7132]*kernel[2]+tmp[7230]*kernel[3]+tmp[7231]*kernel[4]+tmp[7232]*kernel[5]+tmp[7330]*kernel[6]+tmp[7331]*kernel[7]+tmp[7332]*kernel[8];
				ans[7232]<=tmp[7131]*kernel[0]+tmp[7132]*kernel[1]+tmp[7133]*kernel[2]+tmp[7231]*kernel[3]+tmp[7232]*kernel[4]+tmp[7233]*kernel[5]+tmp[7331]*kernel[6]+tmp[7332]*kernel[7]+tmp[7333]*kernel[8];
				ans[7233]<=tmp[7132]*kernel[0]+tmp[7133]*kernel[1]+tmp[7134]*kernel[2]+tmp[7232]*kernel[3]+tmp[7233]*kernel[4]+tmp[7234]*kernel[5]+tmp[7332]*kernel[6]+tmp[7333]*kernel[7]+tmp[7334]*kernel[8];
				ans[7234]<=tmp[7133]*kernel[0]+tmp[7134]*kernel[1]+tmp[7135]*kernel[2]+tmp[7233]*kernel[3]+tmp[7234]*kernel[4]+tmp[7235]*kernel[5]+tmp[7333]*kernel[6]+tmp[7334]*kernel[7]+tmp[7335]*kernel[8];
				ans[7235]<=tmp[7134]*kernel[0]+tmp[7135]*kernel[1]+tmp[7136]*kernel[2]+tmp[7234]*kernel[3]+tmp[7235]*kernel[4]+tmp[7236]*kernel[5]+tmp[7334]*kernel[6]+tmp[7335]*kernel[7]+tmp[7336]*kernel[8];
				ans[7236]<=tmp[7135]*kernel[0]+tmp[7136]*kernel[1]+tmp[7137]*kernel[2]+tmp[7235]*kernel[3]+tmp[7236]*kernel[4]+tmp[7237]*kernel[5]+tmp[7335]*kernel[6]+tmp[7336]*kernel[7]+tmp[7337]*kernel[8];
				ans[7237]<=tmp[7136]*kernel[0]+tmp[7137]*kernel[1]+tmp[7138]*kernel[2]+tmp[7236]*kernel[3]+tmp[7237]*kernel[4]+tmp[7238]*kernel[5]+tmp[7336]*kernel[6]+tmp[7337]*kernel[7]+tmp[7338]*kernel[8];
				ans[7238]<=tmp[7137]*kernel[0]+tmp[7138]*kernel[1]+tmp[7139]*kernel[2]+tmp[7237]*kernel[3]+tmp[7238]*kernel[4]+tmp[7239]*kernel[5]+tmp[7337]*kernel[6]+tmp[7338]*kernel[7]+tmp[7339]*kernel[8];
				ans[7239]<=tmp[7138]*kernel[0]+tmp[7139]*kernel[1]+tmp[7140]*kernel[2]+tmp[7238]*kernel[3]+tmp[7239]*kernel[4]+tmp[7240]*kernel[5]+tmp[7338]*kernel[6]+tmp[7339]*kernel[7]+tmp[7340]*kernel[8];
				ans[7240]<=tmp[7139]*kernel[0]+tmp[7140]*kernel[1]+tmp[7141]*kernel[2]+tmp[7239]*kernel[3]+tmp[7240]*kernel[4]+tmp[7241]*kernel[5]+tmp[7339]*kernel[6]+tmp[7340]*kernel[7]+tmp[7341]*kernel[8];
				ans[7241]<=tmp[7140]*kernel[0]+tmp[7141]*kernel[1]+tmp[7142]*kernel[2]+tmp[7240]*kernel[3]+tmp[7241]*kernel[4]+tmp[7242]*kernel[5]+tmp[7340]*kernel[6]+tmp[7341]*kernel[7]+tmp[7342]*kernel[8];
				ans[7242]<=tmp[7141]*kernel[0]+tmp[7142]*kernel[1]+tmp[7143]*kernel[2]+tmp[7241]*kernel[3]+tmp[7242]*kernel[4]+tmp[7243]*kernel[5]+tmp[7341]*kernel[6]+tmp[7342]*kernel[7]+tmp[7343]*kernel[8];
				ans[7243]<=tmp[7142]*kernel[0]+tmp[7143]*kernel[1]+tmp[7144]*kernel[2]+tmp[7242]*kernel[3]+tmp[7243]*kernel[4]+tmp[7244]*kernel[5]+tmp[7342]*kernel[6]+tmp[7343]*kernel[7]+tmp[7344]*kernel[8];
				ans[7244]<=tmp[7143]*kernel[0]+tmp[7144]*kernel[1]+tmp[7145]*kernel[2]+tmp[7243]*kernel[3]+tmp[7244]*kernel[4]+tmp[7245]*kernel[5]+tmp[7343]*kernel[6]+tmp[7344]*kernel[7]+tmp[7345]*kernel[8];
				ans[7245]<=tmp[7144]*kernel[0]+tmp[7145]*kernel[1]+tmp[7146]*kernel[2]+tmp[7244]*kernel[3]+tmp[7245]*kernel[4]+tmp[7246]*kernel[5]+tmp[7344]*kernel[6]+tmp[7345]*kernel[7]+tmp[7346]*kernel[8];
				ans[7246]<=tmp[7145]*kernel[0]+tmp[7146]*kernel[1]+tmp[7147]*kernel[2]+tmp[7245]*kernel[3]+tmp[7246]*kernel[4]+tmp[7247]*kernel[5]+tmp[7345]*kernel[6]+tmp[7346]*kernel[7]+tmp[7347]*kernel[8];
				ans[7247]<=tmp[7146]*kernel[0]+tmp[7147]*kernel[1]+tmp[7148]*kernel[2]+tmp[7246]*kernel[3]+tmp[7247]*kernel[4]+tmp[7248]*kernel[5]+tmp[7346]*kernel[6]+tmp[7347]*kernel[7]+tmp[7348]*kernel[8];
				ans[7248]<=tmp[7147]*kernel[0]+tmp[7148]*kernel[1]+tmp[7149]*kernel[2]+tmp[7247]*kernel[3]+tmp[7248]*kernel[4]+tmp[7249]*kernel[5]+tmp[7347]*kernel[6]+tmp[7348]*kernel[7]+tmp[7349]*kernel[8];
				ans[7249]<=tmp[7148]*kernel[0]+tmp[7149]*kernel[1]+tmp[7150]*kernel[2]+tmp[7248]*kernel[3]+tmp[7249]*kernel[4]+tmp[7250]*kernel[5]+tmp[7348]*kernel[6]+tmp[7349]*kernel[7]+tmp[7350]*kernel[8];
				ans[7250]<=tmp[7149]*kernel[0]+tmp[7150]*kernel[1]+tmp[7151]*kernel[2]+tmp[7249]*kernel[3]+tmp[7250]*kernel[4]+tmp[7251]*kernel[5]+tmp[7349]*kernel[6]+tmp[7350]*kernel[7]+tmp[7351]*kernel[8];
				ans[7251]<=tmp[7150]*kernel[0]+tmp[7151]*kernel[1]+tmp[7152]*kernel[2]+tmp[7250]*kernel[3]+tmp[7251]*kernel[4]+tmp[7252]*kernel[5]+tmp[7350]*kernel[6]+tmp[7351]*kernel[7]+tmp[7352]*kernel[8];
				ans[7252]<=tmp[7151]*kernel[0]+tmp[7152]*kernel[1]+tmp[7153]*kernel[2]+tmp[7251]*kernel[3]+tmp[7252]*kernel[4]+tmp[7253]*kernel[5]+tmp[7351]*kernel[6]+tmp[7352]*kernel[7]+tmp[7353]*kernel[8];
				ans[7253]<=tmp[7152]*kernel[0]+tmp[7153]*kernel[1]+tmp[7154]*kernel[2]+tmp[7252]*kernel[3]+tmp[7253]*kernel[4]+tmp[7254]*kernel[5]+tmp[7352]*kernel[6]+tmp[7353]*kernel[7]+tmp[7354]*kernel[8];
				ans[7254]<=tmp[7153]*kernel[0]+tmp[7154]*kernel[1]+tmp[7155]*kernel[2]+tmp[7253]*kernel[3]+tmp[7254]*kernel[4]+tmp[7255]*kernel[5]+tmp[7353]*kernel[6]+tmp[7354]*kernel[7]+tmp[7355]*kernel[8];
				ans[7255]<=tmp[7154]*kernel[0]+tmp[7155]*kernel[1]+tmp[7156]*kernel[2]+tmp[7254]*kernel[3]+tmp[7255]*kernel[4]+tmp[7256]*kernel[5]+tmp[7354]*kernel[6]+tmp[7355]*kernel[7]+tmp[7356]*kernel[8];
				ans[7256]<=tmp[7155]*kernel[0]+tmp[7156]*kernel[1]+tmp[7157]*kernel[2]+tmp[7255]*kernel[3]+tmp[7256]*kernel[4]+tmp[7257]*kernel[5]+tmp[7355]*kernel[6]+tmp[7356]*kernel[7]+tmp[7357]*kernel[8];
				ans[7257]<=tmp[7156]*kernel[0]+tmp[7157]*kernel[1]+tmp[7158]*kernel[2]+tmp[7256]*kernel[3]+tmp[7257]*kernel[4]+tmp[7258]*kernel[5]+tmp[7356]*kernel[6]+tmp[7357]*kernel[7]+tmp[7358]*kernel[8];
				ans[7258]<=tmp[7157]*kernel[0]+tmp[7158]*kernel[1]+tmp[7159]*kernel[2]+tmp[7257]*kernel[3]+tmp[7258]*kernel[4]+tmp[7259]*kernel[5]+tmp[7357]*kernel[6]+tmp[7358]*kernel[7]+tmp[7359]*kernel[8];
				ans[7259]<=tmp[7158]*kernel[0]+tmp[7159]*kernel[1]+tmp[7160]*kernel[2]+tmp[7258]*kernel[3]+tmp[7259]*kernel[4]+tmp[7260]*kernel[5]+tmp[7358]*kernel[6]+tmp[7359]*kernel[7]+tmp[7360]*kernel[8];
				ans[7260]<=tmp[7159]*kernel[0]+tmp[7160]*kernel[1]+tmp[7161]*kernel[2]+tmp[7259]*kernel[3]+tmp[7260]*kernel[4]+tmp[7261]*kernel[5]+tmp[7359]*kernel[6]+tmp[7360]*kernel[7]+tmp[7361]*kernel[8];
				ans[7261]<=tmp[7160]*kernel[0]+tmp[7161]*kernel[1]+tmp[7162]*kernel[2]+tmp[7260]*kernel[3]+tmp[7261]*kernel[4]+tmp[7262]*kernel[5]+tmp[7360]*kernel[6]+tmp[7361]*kernel[7]+tmp[7362]*kernel[8];
				ans[7262]<=tmp[7161]*kernel[0]+tmp[7162]*kernel[1]+tmp[7163]*kernel[2]+tmp[7261]*kernel[3]+tmp[7262]*kernel[4]+tmp[7263]*kernel[5]+tmp[7361]*kernel[6]+tmp[7362]*kernel[7]+tmp[7363]*kernel[8];
				ans[7263]<=tmp[7162]*kernel[0]+tmp[7163]*kernel[1]+tmp[7164]*kernel[2]+tmp[7262]*kernel[3]+tmp[7263]*kernel[4]+tmp[7264]*kernel[5]+tmp[7362]*kernel[6]+tmp[7363]*kernel[7]+tmp[7364]*kernel[8];
				ans[7264]<=tmp[7163]*kernel[0]+tmp[7164]*kernel[1]+tmp[7165]*kernel[2]+tmp[7263]*kernel[3]+tmp[7264]*kernel[4]+tmp[7265]*kernel[5]+tmp[7363]*kernel[6]+tmp[7364]*kernel[7]+tmp[7365]*kernel[8];
				ans[7265]<=tmp[7164]*kernel[0]+tmp[7165]*kernel[1]+tmp[7166]*kernel[2]+tmp[7264]*kernel[3]+tmp[7265]*kernel[4]+tmp[7266]*kernel[5]+tmp[7364]*kernel[6]+tmp[7365]*kernel[7]+tmp[7366]*kernel[8];
				ans[7266]<=tmp[7165]*kernel[0]+tmp[7166]*kernel[1]+tmp[7167]*kernel[2]+tmp[7265]*kernel[3]+tmp[7266]*kernel[4]+tmp[7267]*kernel[5]+tmp[7365]*kernel[6]+tmp[7366]*kernel[7]+tmp[7367]*kernel[8];
				ans[7267]<=tmp[7166]*kernel[0]+tmp[7167]*kernel[1]+tmp[7168]*kernel[2]+tmp[7266]*kernel[3]+tmp[7267]*kernel[4]+tmp[7268]*kernel[5]+tmp[7366]*kernel[6]+tmp[7367]*kernel[7]+tmp[7368]*kernel[8];
				ans[7268]<=tmp[7167]*kernel[0]+tmp[7168]*kernel[1]+tmp[7169]*kernel[2]+tmp[7267]*kernel[3]+tmp[7268]*kernel[4]+tmp[7269]*kernel[5]+tmp[7367]*kernel[6]+tmp[7368]*kernel[7]+tmp[7369]*kernel[8];
				ans[7269]<=tmp[7168]*kernel[0]+tmp[7169]*kernel[1]+tmp[7170]*kernel[2]+tmp[7268]*kernel[3]+tmp[7269]*kernel[4]+tmp[7270]*kernel[5]+tmp[7368]*kernel[6]+tmp[7369]*kernel[7]+tmp[7370]*kernel[8];
				ans[7270]<=tmp[7169]*kernel[0]+tmp[7170]*kernel[1]+tmp[7171]*kernel[2]+tmp[7269]*kernel[3]+tmp[7270]*kernel[4]+tmp[7271]*kernel[5]+tmp[7369]*kernel[6]+tmp[7370]*kernel[7]+tmp[7371]*kernel[8];
				ans[7271]<=tmp[7170]*kernel[0]+tmp[7171]*kernel[1]+tmp[7172]*kernel[2]+tmp[7270]*kernel[3]+tmp[7271]*kernel[4]+tmp[7272]*kernel[5]+tmp[7370]*kernel[6]+tmp[7371]*kernel[7]+tmp[7372]*kernel[8];
				ans[7272]<=tmp[7171]*kernel[0]+tmp[7172]*kernel[1]+tmp[7173]*kernel[2]+tmp[7271]*kernel[3]+tmp[7272]*kernel[4]+tmp[7273]*kernel[5]+tmp[7371]*kernel[6]+tmp[7372]*kernel[7]+tmp[7373]*kernel[8];
				ans[7273]<=tmp[7172]*kernel[0]+tmp[7173]*kernel[1]+tmp[7174]*kernel[2]+tmp[7272]*kernel[3]+tmp[7273]*kernel[4]+tmp[7274]*kernel[5]+tmp[7372]*kernel[6]+tmp[7373]*kernel[7]+tmp[7374]*kernel[8];
				ans[7274]<=tmp[7173]*kernel[0]+tmp[7174]*kernel[1]+tmp[7175]*kernel[2]+tmp[7273]*kernel[3]+tmp[7274]*kernel[4]+tmp[7275]*kernel[5]+tmp[7373]*kernel[6]+tmp[7374]*kernel[7]+tmp[7375]*kernel[8];
				ans[7275]<=tmp[7174]*kernel[0]+tmp[7175]*kernel[1]+tmp[7176]*kernel[2]+tmp[7274]*kernel[3]+tmp[7275]*kernel[4]+tmp[7276]*kernel[5]+tmp[7374]*kernel[6]+tmp[7375]*kernel[7]+tmp[7376]*kernel[8];
				ans[7276]<=tmp[7175]*kernel[0]+tmp[7176]*kernel[1]+tmp[7177]*kernel[2]+tmp[7275]*kernel[3]+tmp[7276]*kernel[4]+tmp[7277]*kernel[5]+tmp[7375]*kernel[6]+tmp[7376]*kernel[7]+tmp[7377]*kernel[8];
				ans[7277]<=tmp[7176]*kernel[0]+tmp[7177]*kernel[1]+tmp[7178]*kernel[2]+tmp[7276]*kernel[3]+tmp[7277]*kernel[4]+tmp[7278]*kernel[5]+tmp[7376]*kernel[6]+tmp[7377]*kernel[7]+tmp[7378]*kernel[8];
				ans[7278]<=tmp[7177]*kernel[0]+tmp[7178]*kernel[1]+tmp[7179]*kernel[2]+tmp[7277]*kernel[3]+tmp[7278]*kernel[4]+tmp[7279]*kernel[5]+tmp[7377]*kernel[6]+tmp[7378]*kernel[7]+tmp[7379]*kernel[8];
				ans[7279]<=tmp[7178]*kernel[0]+tmp[7179]*kernel[1]+tmp[7180]*kernel[2]+tmp[7278]*kernel[3]+tmp[7279]*kernel[4]+tmp[7280]*kernel[5]+tmp[7378]*kernel[6]+tmp[7379]*kernel[7]+tmp[7380]*kernel[8];
				ans[7280]<=tmp[7179]*kernel[0]+tmp[7180]*kernel[1]+tmp[7181]*kernel[2]+tmp[7279]*kernel[3]+tmp[7280]*kernel[4]+tmp[7281]*kernel[5]+tmp[7379]*kernel[6]+tmp[7380]*kernel[7]+tmp[7381]*kernel[8];
				ans[7281]<=tmp[7180]*kernel[0]+tmp[7181]*kernel[1]+tmp[7182]*kernel[2]+tmp[7280]*kernel[3]+tmp[7281]*kernel[4]+tmp[7282]*kernel[5]+tmp[7380]*kernel[6]+tmp[7381]*kernel[7]+tmp[7382]*kernel[8];
				ans[7282]<=tmp[7181]*kernel[0]+tmp[7182]*kernel[1]+tmp[7183]*kernel[2]+tmp[7281]*kernel[3]+tmp[7282]*kernel[4]+tmp[7283]*kernel[5]+tmp[7381]*kernel[6]+tmp[7382]*kernel[7]+tmp[7383]*kernel[8];
				ans[7283]<=tmp[7182]*kernel[0]+tmp[7183]*kernel[1]+tmp[7184]*kernel[2]+tmp[7282]*kernel[3]+tmp[7283]*kernel[4]+tmp[7284]*kernel[5]+tmp[7382]*kernel[6]+tmp[7383]*kernel[7]+tmp[7384]*kernel[8];
				ans[7284]<=tmp[7183]*kernel[0]+tmp[7184]*kernel[1]+tmp[7185]*kernel[2]+tmp[7283]*kernel[3]+tmp[7284]*kernel[4]+tmp[7285]*kernel[5]+tmp[7383]*kernel[6]+tmp[7384]*kernel[7]+tmp[7385]*kernel[8];
				ans[7285]<=tmp[7184]*kernel[0]+tmp[7185]*kernel[1]+tmp[7186]*kernel[2]+tmp[7284]*kernel[3]+tmp[7285]*kernel[4]+tmp[7286]*kernel[5]+tmp[7384]*kernel[6]+tmp[7385]*kernel[7]+tmp[7386]*kernel[8];
				ans[7286]<=tmp[7185]*kernel[0]+tmp[7186]*kernel[1]+tmp[7187]*kernel[2]+tmp[7285]*kernel[3]+tmp[7286]*kernel[4]+tmp[7287]*kernel[5]+tmp[7385]*kernel[6]+tmp[7386]*kernel[7]+tmp[7387]*kernel[8];
				ans[7287]<=tmp[7186]*kernel[0]+tmp[7187]*kernel[1]+tmp[7188]*kernel[2]+tmp[7286]*kernel[3]+tmp[7287]*kernel[4]+tmp[7288]*kernel[5]+tmp[7386]*kernel[6]+tmp[7387]*kernel[7]+tmp[7388]*kernel[8];
				ans[7288]<=tmp[7187]*kernel[0]+tmp[7188]*kernel[1]+tmp[7189]*kernel[2]+tmp[7287]*kernel[3]+tmp[7288]*kernel[4]+tmp[7289]*kernel[5]+tmp[7387]*kernel[6]+tmp[7388]*kernel[7]+tmp[7389]*kernel[8];
				ans[7289]<=tmp[7188]*kernel[0]+tmp[7189]*kernel[1]+tmp[7190]*kernel[2]+tmp[7288]*kernel[3]+tmp[7289]*kernel[4]+tmp[7290]*kernel[5]+tmp[7388]*kernel[6]+tmp[7389]*kernel[7]+tmp[7390]*kernel[8];
				ans[7290]<=tmp[7189]*kernel[0]+tmp[7190]*kernel[1]+tmp[7191]*kernel[2]+tmp[7289]*kernel[3]+tmp[7290]*kernel[4]+tmp[7291]*kernel[5]+tmp[7389]*kernel[6]+tmp[7390]*kernel[7]+tmp[7391]*kernel[8];
				ans[7291]<=tmp[7190]*kernel[0]+tmp[7191]*kernel[1]+tmp[7192]*kernel[2]+tmp[7290]*kernel[3]+tmp[7291]*kernel[4]+tmp[7292]*kernel[5]+tmp[7390]*kernel[6]+tmp[7391]*kernel[7]+tmp[7392]*kernel[8];
				ans[7292]<=tmp[7191]*kernel[0]+tmp[7192]*kernel[1]+tmp[7193]*kernel[2]+tmp[7291]*kernel[3]+tmp[7292]*kernel[4]+tmp[7293]*kernel[5]+tmp[7391]*kernel[6]+tmp[7392]*kernel[7]+tmp[7393]*kernel[8];
				ans[7293]<=tmp[7192]*kernel[0]+tmp[7193]*kernel[1]+tmp[7194]*kernel[2]+tmp[7292]*kernel[3]+tmp[7293]*kernel[4]+tmp[7294]*kernel[5]+tmp[7392]*kernel[6]+tmp[7393]*kernel[7]+tmp[7394]*kernel[8];
				ans[7294]<=tmp[7193]*kernel[0]+tmp[7194]*kernel[1]+tmp[7195]*kernel[2]+tmp[7293]*kernel[3]+tmp[7294]*kernel[4]+tmp[7295]*kernel[5]+tmp[7393]*kernel[6]+tmp[7394]*kernel[7]+tmp[7395]*kernel[8];
				ans[7295]<=tmp[7194]*kernel[0]+tmp[7195]*kernel[1]+tmp[7196]*kernel[2]+tmp[7294]*kernel[3]+tmp[7295]*kernel[4]+tmp[7296]*kernel[5]+tmp[7394]*kernel[6]+tmp[7395]*kernel[7]+tmp[7396]*kernel[8];
				ans[7296]<=tmp[7195]*kernel[0]+tmp[7196]*kernel[1]+tmp[7197]*kernel[2]+tmp[7295]*kernel[3]+tmp[7296]*kernel[4]+tmp[7297]*kernel[5]+tmp[7395]*kernel[6]+tmp[7396]*kernel[7]+tmp[7397]*kernel[8];
				ans[7297]<=tmp[7196]*kernel[0]+tmp[7197]*kernel[1]+tmp[7198]*kernel[2]+tmp[7296]*kernel[3]+tmp[7297]*kernel[4]+tmp[7298]*kernel[5]+tmp[7396]*kernel[6]+tmp[7397]*kernel[7]+tmp[7398]*kernel[8];
				ans[7298]<=tmp[7197]*kernel[0]+tmp[7198]*kernel[1]+tmp[7199]*kernel[2]+tmp[7297]*kernel[3]+tmp[7298]*kernel[4]+tmp[7299]*kernel[5]+tmp[7397]*kernel[6]+tmp[7398]*kernel[7]+tmp[7399]*kernel[8];
				ans[7299]<=tmp[7198]*kernel[0]+tmp[7199]*kernel[1]+tmp[7298]*kernel[3]+tmp[7299]*kernel[4]+tmp[7398]*kernel[6]+tmp[7399]*kernel[7];
				ans[7300]<=tmp[7200]*kernel[1]+tmp[7201]*kernel[2]+tmp[7300]*kernel[4]+tmp[7301]*kernel[5]+tmp[7400]*kernel[7]+tmp[7401]*kernel[8];
				ans[7301]<=tmp[7200]*kernel[0]+tmp[7201]*kernel[1]+tmp[7202]*kernel[2]+tmp[7300]*kernel[3]+tmp[7301]*kernel[4]+tmp[7302]*kernel[5]+tmp[7400]*kernel[6]+tmp[7401]*kernel[7]+tmp[7402]*kernel[8];
				ans[7302]<=tmp[7201]*kernel[0]+tmp[7202]*kernel[1]+tmp[7203]*kernel[2]+tmp[7301]*kernel[3]+tmp[7302]*kernel[4]+tmp[7303]*kernel[5]+tmp[7401]*kernel[6]+tmp[7402]*kernel[7]+tmp[7403]*kernel[8];
				ans[7303]<=tmp[7202]*kernel[0]+tmp[7203]*kernel[1]+tmp[7204]*kernel[2]+tmp[7302]*kernel[3]+tmp[7303]*kernel[4]+tmp[7304]*kernel[5]+tmp[7402]*kernel[6]+tmp[7403]*kernel[7]+tmp[7404]*kernel[8];
				ans[7304]<=tmp[7203]*kernel[0]+tmp[7204]*kernel[1]+tmp[7205]*kernel[2]+tmp[7303]*kernel[3]+tmp[7304]*kernel[4]+tmp[7305]*kernel[5]+tmp[7403]*kernel[6]+tmp[7404]*kernel[7]+tmp[7405]*kernel[8];
				ans[7305]<=tmp[7204]*kernel[0]+tmp[7205]*kernel[1]+tmp[7206]*kernel[2]+tmp[7304]*kernel[3]+tmp[7305]*kernel[4]+tmp[7306]*kernel[5]+tmp[7404]*kernel[6]+tmp[7405]*kernel[7]+tmp[7406]*kernel[8];
				ans[7306]<=tmp[7205]*kernel[0]+tmp[7206]*kernel[1]+tmp[7207]*kernel[2]+tmp[7305]*kernel[3]+tmp[7306]*kernel[4]+tmp[7307]*kernel[5]+tmp[7405]*kernel[6]+tmp[7406]*kernel[7]+tmp[7407]*kernel[8];
				ans[7307]<=tmp[7206]*kernel[0]+tmp[7207]*kernel[1]+tmp[7208]*kernel[2]+tmp[7306]*kernel[3]+tmp[7307]*kernel[4]+tmp[7308]*kernel[5]+tmp[7406]*kernel[6]+tmp[7407]*kernel[7]+tmp[7408]*kernel[8];
				ans[7308]<=tmp[7207]*kernel[0]+tmp[7208]*kernel[1]+tmp[7209]*kernel[2]+tmp[7307]*kernel[3]+tmp[7308]*kernel[4]+tmp[7309]*kernel[5]+tmp[7407]*kernel[6]+tmp[7408]*kernel[7]+tmp[7409]*kernel[8];
				ans[7309]<=tmp[7208]*kernel[0]+tmp[7209]*kernel[1]+tmp[7210]*kernel[2]+tmp[7308]*kernel[3]+tmp[7309]*kernel[4]+tmp[7310]*kernel[5]+tmp[7408]*kernel[6]+tmp[7409]*kernel[7]+tmp[7410]*kernel[8];
				ans[7310]<=tmp[7209]*kernel[0]+tmp[7210]*kernel[1]+tmp[7211]*kernel[2]+tmp[7309]*kernel[3]+tmp[7310]*kernel[4]+tmp[7311]*kernel[5]+tmp[7409]*kernel[6]+tmp[7410]*kernel[7]+tmp[7411]*kernel[8];
				ans[7311]<=tmp[7210]*kernel[0]+tmp[7211]*kernel[1]+tmp[7212]*kernel[2]+tmp[7310]*kernel[3]+tmp[7311]*kernel[4]+tmp[7312]*kernel[5]+tmp[7410]*kernel[6]+tmp[7411]*kernel[7]+tmp[7412]*kernel[8];
				ans[7312]<=tmp[7211]*kernel[0]+tmp[7212]*kernel[1]+tmp[7213]*kernel[2]+tmp[7311]*kernel[3]+tmp[7312]*kernel[4]+tmp[7313]*kernel[5]+tmp[7411]*kernel[6]+tmp[7412]*kernel[7]+tmp[7413]*kernel[8];
				ans[7313]<=tmp[7212]*kernel[0]+tmp[7213]*kernel[1]+tmp[7214]*kernel[2]+tmp[7312]*kernel[3]+tmp[7313]*kernel[4]+tmp[7314]*kernel[5]+tmp[7412]*kernel[6]+tmp[7413]*kernel[7]+tmp[7414]*kernel[8];
				ans[7314]<=tmp[7213]*kernel[0]+tmp[7214]*kernel[1]+tmp[7215]*kernel[2]+tmp[7313]*kernel[3]+tmp[7314]*kernel[4]+tmp[7315]*kernel[5]+tmp[7413]*kernel[6]+tmp[7414]*kernel[7]+tmp[7415]*kernel[8];
				ans[7315]<=tmp[7214]*kernel[0]+tmp[7215]*kernel[1]+tmp[7216]*kernel[2]+tmp[7314]*kernel[3]+tmp[7315]*kernel[4]+tmp[7316]*kernel[5]+tmp[7414]*kernel[6]+tmp[7415]*kernel[7]+tmp[7416]*kernel[8];
				ans[7316]<=tmp[7215]*kernel[0]+tmp[7216]*kernel[1]+tmp[7217]*kernel[2]+tmp[7315]*kernel[3]+tmp[7316]*kernel[4]+tmp[7317]*kernel[5]+tmp[7415]*kernel[6]+tmp[7416]*kernel[7]+tmp[7417]*kernel[8];
				ans[7317]<=tmp[7216]*kernel[0]+tmp[7217]*kernel[1]+tmp[7218]*kernel[2]+tmp[7316]*kernel[3]+tmp[7317]*kernel[4]+tmp[7318]*kernel[5]+tmp[7416]*kernel[6]+tmp[7417]*kernel[7]+tmp[7418]*kernel[8];
				ans[7318]<=tmp[7217]*kernel[0]+tmp[7218]*kernel[1]+tmp[7219]*kernel[2]+tmp[7317]*kernel[3]+tmp[7318]*kernel[4]+tmp[7319]*kernel[5]+tmp[7417]*kernel[6]+tmp[7418]*kernel[7]+tmp[7419]*kernel[8];
				ans[7319]<=tmp[7218]*kernel[0]+tmp[7219]*kernel[1]+tmp[7220]*kernel[2]+tmp[7318]*kernel[3]+tmp[7319]*kernel[4]+tmp[7320]*kernel[5]+tmp[7418]*kernel[6]+tmp[7419]*kernel[7]+tmp[7420]*kernel[8];
				ans[7320]<=tmp[7219]*kernel[0]+tmp[7220]*kernel[1]+tmp[7221]*kernel[2]+tmp[7319]*kernel[3]+tmp[7320]*kernel[4]+tmp[7321]*kernel[5]+tmp[7419]*kernel[6]+tmp[7420]*kernel[7]+tmp[7421]*kernel[8];
				ans[7321]<=tmp[7220]*kernel[0]+tmp[7221]*kernel[1]+tmp[7222]*kernel[2]+tmp[7320]*kernel[3]+tmp[7321]*kernel[4]+tmp[7322]*kernel[5]+tmp[7420]*kernel[6]+tmp[7421]*kernel[7]+tmp[7422]*kernel[8];
				ans[7322]<=tmp[7221]*kernel[0]+tmp[7222]*kernel[1]+tmp[7223]*kernel[2]+tmp[7321]*kernel[3]+tmp[7322]*kernel[4]+tmp[7323]*kernel[5]+tmp[7421]*kernel[6]+tmp[7422]*kernel[7]+tmp[7423]*kernel[8];
				ans[7323]<=tmp[7222]*kernel[0]+tmp[7223]*kernel[1]+tmp[7224]*kernel[2]+tmp[7322]*kernel[3]+tmp[7323]*kernel[4]+tmp[7324]*kernel[5]+tmp[7422]*kernel[6]+tmp[7423]*kernel[7]+tmp[7424]*kernel[8];
				ans[7324]<=tmp[7223]*kernel[0]+tmp[7224]*kernel[1]+tmp[7225]*kernel[2]+tmp[7323]*kernel[3]+tmp[7324]*kernel[4]+tmp[7325]*kernel[5]+tmp[7423]*kernel[6]+tmp[7424]*kernel[7]+tmp[7425]*kernel[8];
				ans[7325]<=tmp[7224]*kernel[0]+tmp[7225]*kernel[1]+tmp[7226]*kernel[2]+tmp[7324]*kernel[3]+tmp[7325]*kernel[4]+tmp[7326]*kernel[5]+tmp[7424]*kernel[6]+tmp[7425]*kernel[7]+tmp[7426]*kernel[8];
				ans[7326]<=tmp[7225]*kernel[0]+tmp[7226]*kernel[1]+tmp[7227]*kernel[2]+tmp[7325]*kernel[3]+tmp[7326]*kernel[4]+tmp[7327]*kernel[5]+tmp[7425]*kernel[6]+tmp[7426]*kernel[7]+tmp[7427]*kernel[8];
				ans[7327]<=tmp[7226]*kernel[0]+tmp[7227]*kernel[1]+tmp[7228]*kernel[2]+tmp[7326]*kernel[3]+tmp[7327]*kernel[4]+tmp[7328]*kernel[5]+tmp[7426]*kernel[6]+tmp[7427]*kernel[7]+tmp[7428]*kernel[8];
				ans[7328]<=tmp[7227]*kernel[0]+tmp[7228]*kernel[1]+tmp[7229]*kernel[2]+tmp[7327]*kernel[3]+tmp[7328]*kernel[4]+tmp[7329]*kernel[5]+tmp[7427]*kernel[6]+tmp[7428]*kernel[7]+tmp[7429]*kernel[8];
				ans[7329]<=tmp[7228]*kernel[0]+tmp[7229]*kernel[1]+tmp[7230]*kernel[2]+tmp[7328]*kernel[3]+tmp[7329]*kernel[4]+tmp[7330]*kernel[5]+tmp[7428]*kernel[6]+tmp[7429]*kernel[7]+tmp[7430]*kernel[8];
				ans[7330]<=tmp[7229]*kernel[0]+tmp[7230]*kernel[1]+tmp[7231]*kernel[2]+tmp[7329]*kernel[3]+tmp[7330]*kernel[4]+tmp[7331]*kernel[5]+tmp[7429]*kernel[6]+tmp[7430]*kernel[7]+tmp[7431]*kernel[8];
				ans[7331]<=tmp[7230]*kernel[0]+tmp[7231]*kernel[1]+tmp[7232]*kernel[2]+tmp[7330]*kernel[3]+tmp[7331]*kernel[4]+tmp[7332]*kernel[5]+tmp[7430]*kernel[6]+tmp[7431]*kernel[7]+tmp[7432]*kernel[8];
				ans[7332]<=tmp[7231]*kernel[0]+tmp[7232]*kernel[1]+tmp[7233]*kernel[2]+tmp[7331]*kernel[3]+tmp[7332]*kernel[4]+tmp[7333]*kernel[5]+tmp[7431]*kernel[6]+tmp[7432]*kernel[7]+tmp[7433]*kernel[8];
				ans[7333]<=tmp[7232]*kernel[0]+tmp[7233]*kernel[1]+tmp[7234]*kernel[2]+tmp[7332]*kernel[3]+tmp[7333]*kernel[4]+tmp[7334]*kernel[5]+tmp[7432]*kernel[6]+tmp[7433]*kernel[7]+tmp[7434]*kernel[8];
				ans[7334]<=tmp[7233]*kernel[0]+tmp[7234]*kernel[1]+tmp[7235]*kernel[2]+tmp[7333]*kernel[3]+tmp[7334]*kernel[4]+tmp[7335]*kernel[5]+tmp[7433]*kernel[6]+tmp[7434]*kernel[7]+tmp[7435]*kernel[8];
				ans[7335]<=tmp[7234]*kernel[0]+tmp[7235]*kernel[1]+tmp[7236]*kernel[2]+tmp[7334]*kernel[3]+tmp[7335]*kernel[4]+tmp[7336]*kernel[5]+tmp[7434]*kernel[6]+tmp[7435]*kernel[7]+tmp[7436]*kernel[8];
				ans[7336]<=tmp[7235]*kernel[0]+tmp[7236]*kernel[1]+tmp[7237]*kernel[2]+tmp[7335]*kernel[3]+tmp[7336]*kernel[4]+tmp[7337]*kernel[5]+tmp[7435]*kernel[6]+tmp[7436]*kernel[7]+tmp[7437]*kernel[8];
				ans[7337]<=tmp[7236]*kernel[0]+tmp[7237]*kernel[1]+tmp[7238]*kernel[2]+tmp[7336]*kernel[3]+tmp[7337]*kernel[4]+tmp[7338]*kernel[5]+tmp[7436]*kernel[6]+tmp[7437]*kernel[7]+tmp[7438]*kernel[8];
				ans[7338]<=tmp[7237]*kernel[0]+tmp[7238]*kernel[1]+tmp[7239]*kernel[2]+tmp[7337]*kernel[3]+tmp[7338]*kernel[4]+tmp[7339]*kernel[5]+tmp[7437]*kernel[6]+tmp[7438]*kernel[7]+tmp[7439]*kernel[8];
				ans[7339]<=tmp[7238]*kernel[0]+tmp[7239]*kernel[1]+tmp[7240]*kernel[2]+tmp[7338]*kernel[3]+tmp[7339]*kernel[4]+tmp[7340]*kernel[5]+tmp[7438]*kernel[6]+tmp[7439]*kernel[7]+tmp[7440]*kernel[8];
				ans[7340]<=tmp[7239]*kernel[0]+tmp[7240]*kernel[1]+tmp[7241]*kernel[2]+tmp[7339]*kernel[3]+tmp[7340]*kernel[4]+tmp[7341]*kernel[5]+tmp[7439]*kernel[6]+tmp[7440]*kernel[7]+tmp[7441]*kernel[8];
				ans[7341]<=tmp[7240]*kernel[0]+tmp[7241]*kernel[1]+tmp[7242]*kernel[2]+tmp[7340]*kernel[3]+tmp[7341]*kernel[4]+tmp[7342]*kernel[5]+tmp[7440]*kernel[6]+tmp[7441]*kernel[7]+tmp[7442]*kernel[8];
				ans[7342]<=tmp[7241]*kernel[0]+tmp[7242]*kernel[1]+tmp[7243]*kernel[2]+tmp[7341]*kernel[3]+tmp[7342]*kernel[4]+tmp[7343]*kernel[5]+tmp[7441]*kernel[6]+tmp[7442]*kernel[7]+tmp[7443]*kernel[8];
				ans[7343]<=tmp[7242]*kernel[0]+tmp[7243]*kernel[1]+tmp[7244]*kernel[2]+tmp[7342]*kernel[3]+tmp[7343]*kernel[4]+tmp[7344]*kernel[5]+tmp[7442]*kernel[6]+tmp[7443]*kernel[7]+tmp[7444]*kernel[8];
				ans[7344]<=tmp[7243]*kernel[0]+tmp[7244]*kernel[1]+tmp[7245]*kernel[2]+tmp[7343]*kernel[3]+tmp[7344]*kernel[4]+tmp[7345]*kernel[5]+tmp[7443]*kernel[6]+tmp[7444]*kernel[7]+tmp[7445]*kernel[8];
				ans[7345]<=tmp[7244]*kernel[0]+tmp[7245]*kernel[1]+tmp[7246]*kernel[2]+tmp[7344]*kernel[3]+tmp[7345]*kernel[4]+tmp[7346]*kernel[5]+tmp[7444]*kernel[6]+tmp[7445]*kernel[7]+tmp[7446]*kernel[8];
				ans[7346]<=tmp[7245]*kernel[0]+tmp[7246]*kernel[1]+tmp[7247]*kernel[2]+tmp[7345]*kernel[3]+tmp[7346]*kernel[4]+tmp[7347]*kernel[5]+tmp[7445]*kernel[6]+tmp[7446]*kernel[7]+tmp[7447]*kernel[8];
				ans[7347]<=tmp[7246]*kernel[0]+tmp[7247]*kernel[1]+tmp[7248]*kernel[2]+tmp[7346]*kernel[3]+tmp[7347]*kernel[4]+tmp[7348]*kernel[5]+tmp[7446]*kernel[6]+tmp[7447]*kernel[7]+tmp[7448]*kernel[8];
				ans[7348]<=tmp[7247]*kernel[0]+tmp[7248]*kernel[1]+tmp[7249]*kernel[2]+tmp[7347]*kernel[3]+tmp[7348]*kernel[4]+tmp[7349]*kernel[5]+tmp[7447]*kernel[6]+tmp[7448]*kernel[7]+tmp[7449]*kernel[8];
				ans[7349]<=tmp[7248]*kernel[0]+tmp[7249]*kernel[1]+tmp[7250]*kernel[2]+tmp[7348]*kernel[3]+tmp[7349]*kernel[4]+tmp[7350]*kernel[5]+tmp[7448]*kernel[6]+tmp[7449]*kernel[7]+tmp[7450]*kernel[8];
				ans[7350]<=tmp[7249]*kernel[0]+tmp[7250]*kernel[1]+tmp[7251]*kernel[2]+tmp[7349]*kernel[3]+tmp[7350]*kernel[4]+tmp[7351]*kernel[5]+tmp[7449]*kernel[6]+tmp[7450]*kernel[7]+tmp[7451]*kernel[8];
				ans[7351]<=tmp[7250]*kernel[0]+tmp[7251]*kernel[1]+tmp[7252]*kernel[2]+tmp[7350]*kernel[3]+tmp[7351]*kernel[4]+tmp[7352]*kernel[5]+tmp[7450]*kernel[6]+tmp[7451]*kernel[7]+tmp[7452]*kernel[8];
				ans[7352]<=tmp[7251]*kernel[0]+tmp[7252]*kernel[1]+tmp[7253]*kernel[2]+tmp[7351]*kernel[3]+tmp[7352]*kernel[4]+tmp[7353]*kernel[5]+tmp[7451]*kernel[6]+tmp[7452]*kernel[7]+tmp[7453]*kernel[8];
				ans[7353]<=tmp[7252]*kernel[0]+tmp[7253]*kernel[1]+tmp[7254]*kernel[2]+tmp[7352]*kernel[3]+tmp[7353]*kernel[4]+tmp[7354]*kernel[5]+tmp[7452]*kernel[6]+tmp[7453]*kernel[7]+tmp[7454]*kernel[8];
				ans[7354]<=tmp[7253]*kernel[0]+tmp[7254]*kernel[1]+tmp[7255]*kernel[2]+tmp[7353]*kernel[3]+tmp[7354]*kernel[4]+tmp[7355]*kernel[5]+tmp[7453]*kernel[6]+tmp[7454]*kernel[7]+tmp[7455]*kernel[8];
				ans[7355]<=tmp[7254]*kernel[0]+tmp[7255]*kernel[1]+tmp[7256]*kernel[2]+tmp[7354]*kernel[3]+tmp[7355]*kernel[4]+tmp[7356]*kernel[5]+tmp[7454]*kernel[6]+tmp[7455]*kernel[7]+tmp[7456]*kernel[8];
				ans[7356]<=tmp[7255]*kernel[0]+tmp[7256]*kernel[1]+tmp[7257]*kernel[2]+tmp[7355]*kernel[3]+tmp[7356]*kernel[4]+tmp[7357]*kernel[5]+tmp[7455]*kernel[6]+tmp[7456]*kernel[7]+tmp[7457]*kernel[8];
				ans[7357]<=tmp[7256]*kernel[0]+tmp[7257]*kernel[1]+tmp[7258]*kernel[2]+tmp[7356]*kernel[3]+tmp[7357]*kernel[4]+tmp[7358]*kernel[5]+tmp[7456]*kernel[6]+tmp[7457]*kernel[7]+tmp[7458]*kernel[8];
				ans[7358]<=tmp[7257]*kernel[0]+tmp[7258]*kernel[1]+tmp[7259]*kernel[2]+tmp[7357]*kernel[3]+tmp[7358]*kernel[4]+tmp[7359]*kernel[5]+tmp[7457]*kernel[6]+tmp[7458]*kernel[7]+tmp[7459]*kernel[8];
				ans[7359]<=tmp[7258]*kernel[0]+tmp[7259]*kernel[1]+tmp[7260]*kernel[2]+tmp[7358]*kernel[3]+tmp[7359]*kernel[4]+tmp[7360]*kernel[5]+tmp[7458]*kernel[6]+tmp[7459]*kernel[7]+tmp[7460]*kernel[8];
				ans[7360]<=tmp[7259]*kernel[0]+tmp[7260]*kernel[1]+tmp[7261]*kernel[2]+tmp[7359]*kernel[3]+tmp[7360]*kernel[4]+tmp[7361]*kernel[5]+tmp[7459]*kernel[6]+tmp[7460]*kernel[7]+tmp[7461]*kernel[8];
				ans[7361]<=tmp[7260]*kernel[0]+tmp[7261]*kernel[1]+tmp[7262]*kernel[2]+tmp[7360]*kernel[3]+tmp[7361]*kernel[4]+tmp[7362]*kernel[5]+tmp[7460]*kernel[6]+tmp[7461]*kernel[7]+tmp[7462]*kernel[8];
				ans[7362]<=tmp[7261]*kernel[0]+tmp[7262]*kernel[1]+tmp[7263]*kernel[2]+tmp[7361]*kernel[3]+tmp[7362]*kernel[4]+tmp[7363]*kernel[5]+tmp[7461]*kernel[6]+tmp[7462]*kernel[7]+tmp[7463]*kernel[8];
				ans[7363]<=tmp[7262]*kernel[0]+tmp[7263]*kernel[1]+tmp[7264]*kernel[2]+tmp[7362]*kernel[3]+tmp[7363]*kernel[4]+tmp[7364]*kernel[5]+tmp[7462]*kernel[6]+tmp[7463]*kernel[7]+tmp[7464]*kernel[8];
				ans[7364]<=tmp[7263]*kernel[0]+tmp[7264]*kernel[1]+tmp[7265]*kernel[2]+tmp[7363]*kernel[3]+tmp[7364]*kernel[4]+tmp[7365]*kernel[5]+tmp[7463]*kernel[6]+tmp[7464]*kernel[7]+tmp[7465]*kernel[8];
				ans[7365]<=tmp[7264]*kernel[0]+tmp[7265]*kernel[1]+tmp[7266]*kernel[2]+tmp[7364]*kernel[3]+tmp[7365]*kernel[4]+tmp[7366]*kernel[5]+tmp[7464]*kernel[6]+tmp[7465]*kernel[7]+tmp[7466]*kernel[8];
				ans[7366]<=tmp[7265]*kernel[0]+tmp[7266]*kernel[1]+tmp[7267]*kernel[2]+tmp[7365]*kernel[3]+tmp[7366]*kernel[4]+tmp[7367]*kernel[5]+tmp[7465]*kernel[6]+tmp[7466]*kernel[7]+tmp[7467]*kernel[8];
				ans[7367]<=tmp[7266]*kernel[0]+tmp[7267]*kernel[1]+tmp[7268]*kernel[2]+tmp[7366]*kernel[3]+tmp[7367]*kernel[4]+tmp[7368]*kernel[5]+tmp[7466]*kernel[6]+tmp[7467]*kernel[7]+tmp[7468]*kernel[8];
				ans[7368]<=tmp[7267]*kernel[0]+tmp[7268]*kernel[1]+tmp[7269]*kernel[2]+tmp[7367]*kernel[3]+tmp[7368]*kernel[4]+tmp[7369]*kernel[5]+tmp[7467]*kernel[6]+tmp[7468]*kernel[7]+tmp[7469]*kernel[8];
				ans[7369]<=tmp[7268]*kernel[0]+tmp[7269]*kernel[1]+tmp[7270]*kernel[2]+tmp[7368]*kernel[3]+tmp[7369]*kernel[4]+tmp[7370]*kernel[5]+tmp[7468]*kernel[6]+tmp[7469]*kernel[7]+tmp[7470]*kernel[8];
				ans[7370]<=tmp[7269]*kernel[0]+tmp[7270]*kernel[1]+tmp[7271]*kernel[2]+tmp[7369]*kernel[3]+tmp[7370]*kernel[4]+tmp[7371]*kernel[5]+tmp[7469]*kernel[6]+tmp[7470]*kernel[7]+tmp[7471]*kernel[8];
				ans[7371]<=tmp[7270]*kernel[0]+tmp[7271]*kernel[1]+tmp[7272]*kernel[2]+tmp[7370]*kernel[3]+tmp[7371]*kernel[4]+tmp[7372]*kernel[5]+tmp[7470]*kernel[6]+tmp[7471]*kernel[7]+tmp[7472]*kernel[8];
				ans[7372]<=tmp[7271]*kernel[0]+tmp[7272]*kernel[1]+tmp[7273]*kernel[2]+tmp[7371]*kernel[3]+tmp[7372]*kernel[4]+tmp[7373]*kernel[5]+tmp[7471]*kernel[6]+tmp[7472]*kernel[7]+tmp[7473]*kernel[8];
				ans[7373]<=tmp[7272]*kernel[0]+tmp[7273]*kernel[1]+tmp[7274]*kernel[2]+tmp[7372]*kernel[3]+tmp[7373]*kernel[4]+tmp[7374]*kernel[5]+tmp[7472]*kernel[6]+tmp[7473]*kernel[7]+tmp[7474]*kernel[8];
				ans[7374]<=tmp[7273]*kernel[0]+tmp[7274]*kernel[1]+tmp[7275]*kernel[2]+tmp[7373]*kernel[3]+tmp[7374]*kernel[4]+tmp[7375]*kernel[5]+tmp[7473]*kernel[6]+tmp[7474]*kernel[7]+tmp[7475]*kernel[8];
				ans[7375]<=tmp[7274]*kernel[0]+tmp[7275]*kernel[1]+tmp[7276]*kernel[2]+tmp[7374]*kernel[3]+tmp[7375]*kernel[4]+tmp[7376]*kernel[5]+tmp[7474]*kernel[6]+tmp[7475]*kernel[7]+tmp[7476]*kernel[8];
				ans[7376]<=tmp[7275]*kernel[0]+tmp[7276]*kernel[1]+tmp[7277]*kernel[2]+tmp[7375]*kernel[3]+tmp[7376]*kernel[4]+tmp[7377]*kernel[5]+tmp[7475]*kernel[6]+tmp[7476]*kernel[7]+tmp[7477]*kernel[8];
				ans[7377]<=tmp[7276]*kernel[0]+tmp[7277]*kernel[1]+tmp[7278]*kernel[2]+tmp[7376]*kernel[3]+tmp[7377]*kernel[4]+tmp[7378]*kernel[5]+tmp[7476]*kernel[6]+tmp[7477]*kernel[7]+tmp[7478]*kernel[8];
				ans[7378]<=tmp[7277]*kernel[0]+tmp[7278]*kernel[1]+tmp[7279]*kernel[2]+tmp[7377]*kernel[3]+tmp[7378]*kernel[4]+tmp[7379]*kernel[5]+tmp[7477]*kernel[6]+tmp[7478]*kernel[7]+tmp[7479]*kernel[8];
				ans[7379]<=tmp[7278]*kernel[0]+tmp[7279]*kernel[1]+tmp[7280]*kernel[2]+tmp[7378]*kernel[3]+tmp[7379]*kernel[4]+tmp[7380]*kernel[5]+tmp[7478]*kernel[6]+tmp[7479]*kernel[7]+tmp[7480]*kernel[8];
				ans[7380]<=tmp[7279]*kernel[0]+tmp[7280]*kernel[1]+tmp[7281]*kernel[2]+tmp[7379]*kernel[3]+tmp[7380]*kernel[4]+tmp[7381]*kernel[5]+tmp[7479]*kernel[6]+tmp[7480]*kernel[7]+tmp[7481]*kernel[8];
				ans[7381]<=tmp[7280]*kernel[0]+tmp[7281]*kernel[1]+tmp[7282]*kernel[2]+tmp[7380]*kernel[3]+tmp[7381]*kernel[4]+tmp[7382]*kernel[5]+tmp[7480]*kernel[6]+tmp[7481]*kernel[7]+tmp[7482]*kernel[8];
				ans[7382]<=tmp[7281]*kernel[0]+tmp[7282]*kernel[1]+tmp[7283]*kernel[2]+tmp[7381]*kernel[3]+tmp[7382]*kernel[4]+tmp[7383]*kernel[5]+tmp[7481]*kernel[6]+tmp[7482]*kernel[7]+tmp[7483]*kernel[8];
				ans[7383]<=tmp[7282]*kernel[0]+tmp[7283]*kernel[1]+tmp[7284]*kernel[2]+tmp[7382]*kernel[3]+tmp[7383]*kernel[4]+tmp[7384]*kernel[5]+tmp[7482]*kernel[6]+tmp[7483]*kernel[7]+tmp[7484]*kernel[8];
				ans[7384]<=tmp[7283]*kernel[0]+tmp[7284]*kernel[1]+tmp[7285]*kernel[2]+tmp[7383]*kernel[3]+tmp[7384]*kernel[4]+tmp[7385]*kernel[5]+tmp[7483]*kernel[6]+tmp[7484]*kernel[7]+tmp[7485]*kernel[8];
				ans[7385]<=tmp[7284]*kernel[0]+tmp[7285]*kernel[1]+tmp[7286]*kernel[2]+tmp[7384]*kernel[3]+tmp[7385]*kernel[4]+tmp[7386]*kernel[5]+tmp[7484]*kernel[6]+tmp[7485]*kernel[7]+tmp[7486]*kernel[8];
				ans[7386]<=tmp[7285]*kernel[0]+tmp[7286]*kernel[1]+tmp[7287]*kernel[2]+tmp[7385]*kernel[3]+tmp[7386]*kernel[4]+tmp[7387]*kernel[5]+tmp[7485]*kernel[6]+tmp[7486]*kernel[7]+tmp[7487]*kernel[8];
				ans[7387]<=tmp[7286]*kernel[0]+tmp[7287]*kernel[1]+tmp[7288]*kernel[2]+tmp[7386]*kernel[3]+tmp[7387]*kernel[4]+tmp[7388]*kernel[5]+tmp[7486]*kernel[6]+tmp[7487]*kernel[7]+tmp[7488]*kernel[8];
				ans[7388]<=tmp[7287]*kernel[0]+tmp[7288]*kernel[1]+tmp[7289]*kernel[2]+tmp[7387]*kernel[3]+tmp[7388]*kernel[4]+tmp[7389]*kernel[5]+tmp[7487]*kernel[6]+tmp[7488]*kernel[7]+tmp[7489]*kernel[8];
				ans[7389]<=tmp[7288]*kernel[0]+tmp[7289]*kernel[1]+tmp[7290]*kernel[2]+tmp[7388]*kernel[3]+tmp[7389]*kernel[4]+tmp[7390]*kernel[5]+tmp[7488]*kernel[6]+tmp[7489]*kernel[7]+tmp[7490]*kernel[8];
				ans[7390]<=tmp[7289]*kernel[0]+tmp[7290]*kernel[1]+tmp[7291]*kernel[2]+tmp[7389]*kernel[3]+tmp[7390]*kernel[4]+tmp[7391]*kernel[5]+tmp[7489]*kernel[6]+tmp[7490]*kernel[7]+tmp[7491]*kernel[8];
				ans[7391]<=tmp[7290]*kernel[0]+tmp[7291]*kernel[1]+tmp[7292]*kernel[2]+tmp[7390]*kernel[3]+tmp[7391]*kernel[4]+tmp[7392]*kernel[5]+tmp[7490]*kernel[6]+tmp[7491]*kernel[7]+tmp[7492]*kernel[8];
				ans[7392]<=tmp[7291]*kernel[0]+tmp[7292]*kernel[1]+tmp[7293]*kernel[2]+tmp[7391]*kernel[3]+tmp[7392]*kernel[4]+tmp[7393]*kernel[5]+tmp[7491]*kernel[6]+tmp[7492]*kernel[7]+tmp[7493]*kernel[8];
				ans[7393]<=tmp[7292]*kernel[0]+tmp[7293]*kernel[1]+tmp[7294]*kernel[2]+tmp[7392]*kernel[3]+tmp[7393]*kernel[4]+tmp[7394]*kernel[5]+tmp[7492]*kernel[6]+tmp[7493]*kernel[7]+tmp[7494]*kernel[8];
				ans[7394]<=tmp[7293]*kernel[0]+tmp[7294]*kernel[1]+tmp[7295]*kernel[2]+tmp[7393]*kernel[3]+tmp[7394]*kernel[4]+tmp[7395]*kernel[5]+tmp[7493]*kernel[6]+tmp[7494]*kernel[7]+tmp[7495]*kernel[8];
				ans[7395]<=tmp[7294]*kernel[0]+tmp[7295]*kernel[1]+tmp[7296]*kernel[2]+tmp[7394]*kernel[3]+tmp[7395]*kernel[4]+tmp[7396]*kernel[5]+tmp[7494]*kernel[6]+tmp[7495]*kernel[7]+tmp[7496]*kernel[8];
				ans[7396]<=tmp[7295]*kernel[0]+tmp[7296]*kernel[1]+tmp[7297]*kernel[2]+tmp[7395]*kernel[3]+tmp[7396]*kernel[4]+tmp[7397]*kernel[5]+tmp[7495]*kernel[6]+tmp[7496]*kernel[7]+tmp[7497]*kernel[8];
				ans[7397]<=tmp[7296]*kernel[0]+tmp[7297]*kernel[1]+tmp[7298]*kernel[2]+tmp[7396]*kernel[3]+tmp[7397]*kernel[4]+tmp[7398]*kernel[5]+tmp[7496]*kernel[6]+tmp[7497]*kernel[7]+tmp[7498]*kernel[8];
				ans[7398]<=tmp[7297]*kernel[0]+tmp[7298]*kernel[1]+tmp[7299]*kernel[2]+tmp[7397]*kernel[3]+tmp[7398]*kernel[4]+tmp[7399]*kernel[5]+tmp[7497]*kernel[6]+tmp[7498]*kernel[7]+tmp[7499]*kernel[8];
				ans[7399]<=tmp[7298]*kernel[0]+tmp[7299]*kernel[1]+tmp[7398]*kernel[3]+tmp[7399]*kernel[4]+tmp[7498]*kernel[6]+tmp[7499]*kernel[7];
				ans[7400]<=tmp[7300]*kernel[1]+tmp[7301]*kernel[2]+tmp[7400]*kernel[4]+tmp[7401]*kernel[5]+tmp[7500]*kernel[7]+tmp[7501]*kernel[8];
				ans[7401]<=tmp[7300]*kernel[0]+tmp[7301]*kernel[1]+tmp[7302]*kernel[2]+tmp[7400]*kernel[3]+tmp[7401]*kernel[4]+tmp[7402]*kernel[5]+tmp[7500]*kernel[6]+tmp[7501]*kernel[7]+tmp[7502]*kernel[8];
				ans[7402]<=tmp[7301]*kernel[0]+tmp[7302]*kernel[1]+tmp[7303]*kernel[2]+tmp[7401]*kernel[3]+tmp[7402]*kernel[4]+tmp[7403]*kernel[5]+tmp[7501]*kernel[6]+tmp[7502]*kernel[7]+tmp[7503]*kernel[8];
				ans[7403]<=tmp[7302]*kernel[0]+tmp[7303]*kernel[1]+tmp[7304]*kernel[2]+tmp[7402]*kernel[3]+tmp[7403]*kernel[4]+tmp[7404]*kernel[5]+tmp[7502]*kernel[6]+tmp[7503]*kernel[7]+tmp[7504]*kernel[8];
				ans[7404]<=tmp[7303]*kernel[0]+tmp[7304]*kernel[1]+tmp[7305]*kernel[2]+tmp[7403]*kernel[3]+tmp[7404]*kernel[4]+tmp[7405]*kernel[5]+tmp[7503]*kernel[6]+tmp[7504]*kernel[7]+tmp[7505]*kernel[8];
				ans[7405]<=tmp[7304]*kernel[0]+tmp[7305]*kernel[1]+tmp[7306]*kernel[2]+tmp[7404]*kernel[3]+tmp[7405]*kernel[4]+tmp[7406]*kernel[5]+tmp[7504]*kernel[6]+tmp[7505]*kernel[7]+tmp[7506]*kernel[8];
				ans[7406]<=tmp[7305]*kernel[0]+tmp[7306]*kernel[1]+tmp[7307]*kernel[2]+tmp[7405]*kernel[3]+tmp[7406]*kernel[4]+tmp[7407]*kernel[5]+tmp[7505]*kernel[6]+tmp[7506]*kernel[7]+tmp[7507]*kernel[8];
				ans[7407]<=tmp[7306]*kernel[0]+tmp[7307]*kernel[1]+tmp[7308]*kernel[2]+tmp[7406]*kernel[3]+tmp[7407]*kernel[4]+tmp[7408]*kernel[5]+tmp[7506]*kernel[6]+tmp[7507]*kernel[7]+tmp[7508]*kernel[8];
				ans[7408]<=tmp[7307]*kernel[0]+tmp[7308]*kernel[1]+tmp[7309]*kernel[2]+tmp[7407]*kernel[3]+tmp[7408]*kernel[4]+tmp[7409]*kernel[5]+tmp[7507]*kernel[6]+tmp[7508]*kernel[7]+tmp[7509]*kernel[8];
				ans[7409]<=tmp[7308]*kernel[0]+tmp[7309]*kernel[1]+tmp[7310]*kernel[2]+tmp[7408]*kernel[3]+tmp[7409]*kernel[4]+tmp[7410]*kernel[5]+tmp[7508]*kernel[6]+tmp[7509]*kernel[7]+tmp[7510]*kernel[8];
				ans[7410]<=tmp[7309]*kernel[0]+tmp[7310]*kernel[1]+tmp[7311]*kernel[2]+tmp[7409]*kernel[3]+tmp[7410]*kernel[4]+tmp[7411]*kernel[5]+tmp[7509]*kernel[6]+tmp[7510]*kernel[7]+tmp[7511]*kernel[8];
				ans[7411]<=tmp[7310]*kernel[0]+tmp[7311]*kernel[1]+tmp[7312]*kernel[2]+tmp[7410]*kernel[3]+tmp[7411]*kernel[4]+tmp[7412]*kernel[5]+tmp[7510]*kernel[6]+tmp[7511]*kernel[7]+tmp[7512]*kernel[8];
				ans[7412]<=tmp[7311]*kernel[0]+tmp[7312]*kernel[1]+tmp[7313]*kernel[2]+tmp[7411]*kernel[3]+tmp[7412]*kernel[4]+tmp[7413]*kernel[5]+tmp[7511]*kernel[6]+tmp[7512]*kernel[7]+tmp[7513]*kernel[8];
				ans[7413]<=tmp[7312]*kernel[0]+tmp[7313]*kernel[1]+tmp[7314]*kernel[2]+tmp[7412]*kernel[3]+tmp[7413]*kernel[4]+tmp[7414]*kernel[5]+tmp[7512]*kernel[6]+tmp[7513]*kernel[7]+tmp[7514]*kernel[8];
				ans[7414]<=tmp[7313]*kernel[0]+tmp[7314]*kernel[1]+tmp[7315]*kernel[2]+tmp[7413]*kernel[3]+tmp[7414]*kernel[4]+tmp[7415]*kernel[5]+tmp[7513]*kernel[6]+tmp[7514]*kernel[7]+tmp[7515]*kernel[8];
				ans[7415]<=tmp[7314]*kernel[0]+tmp[7315]*kernel[1]+tmp[7316]*kernel[2]+tmp[7414]*kernel[3]+tmp[7415]*kernel[4]+tmp[7416]*kernel[5]+tmp[7514]*kernel[6]+tmp[7515]*kernel[7]+tmp[7516]*kernel[8];
				ans[7416]<=tmp[7315]*kernel[0]+tmp[7316]*kernel[1]+tmp[7317]*kernel[2]+tmp[7415]*kernel[3]+tmp[7416]*kernel[4]+tmp[7417]*kernel[5]+tmp[7515]*kernel[6]+tmp[7516]*kernel[7]+tmp[7517]*kernel[8];
				ans[7417]<=tmp[7316]*kernel[0]+tmp[7317]*kernel[1]+tmp[7318]*kernel[2]+tmp[7416]*kernel[3]+tmp[7417]*kernel[4]+tmp[7418]*kernel[5]+tmp[7516]*kernel[6]+tmp[7517]*kernel[7]+tmp[7518]*kernel[8];
				ans[7418]<=tmp[7317]*kernel[0]+tmp[7318]*kernel[1]+tmp[7319]*kernel[2]+tmp[7417]*kernel[3]+tmp[7418]*kernel[4]+tmp[7419]*kernel[5]+tmp[7517]*kernel[6]+tmp[7518]*kernel[7]+tmp[7519]*kernel[8];
				ans[7419]<=tmp[7318]*kernel[0]+tmp[7319]*kernel[1]+tmp[7320]*kernel[2]+tmp[7418]*kernel[3]+tmp[7419]*kernel[4]+tmp[7420]*kernel[5]+tmp[7518]*kernel[6]+tmp[7519]*kernel[7]+tmp[7520]*kernel[8];
				ans[7420]<=tmp[7319]*kernel[0]+tmp[7320]*kernel[1]+tmp[7321]*kernel[2]+tmp[7419]*kernel[3]+tmp[7420]*kernel[4]+tmp[7421]*kernel[5]+tmp[7519]*kernel[6]+tmp[7520]*kernel[7]+tmp[7521]*kernel[8];
				ans[7421]<=tmp[7320]*kernel[0]+tmp[7321]*kernel[1]+tmp[7322]*kernel[2]+tmp[7420]*kernel[3]+tmp[7421]*kernel[4]+tmp[7422]*kernel[5]+tmp[7520]*kernel[6]+tmp[7521]*kernel[7]+tmp[7522]*kernel[8];
				ans[7422]<=tmp[7321]*kernel[0]+tmp[7322]*kernel[1]+tmp[7323]*kernel[2]+tmp[7421]*kernel[3]+tmp[7422]*kernel[4]+tmp[7423]*kernel[5]+tmp[7521]*kernel[6]+tmp[7522]*kernel[7]+tmp[7523]*kernel[8];
				ans[7423]<=tmp[7322]*kernel[0]+tmp[7323]*kernel[1]+tmp[7324]*kernel[2]+tmp[7422]*kernel[3]+tmp[7423]*kernel[4]+tmp[7424]*kernel[5]+tmp[7522]*kernel[6]+tmp[7523]*kernel[7]+tmp[7524]*kernel[8];
				ans[7424]<=tmp[7323]*kernel[0]+tmp[7324]*kernel[1]+tmp[7325]*kernel[2]+tmp[7423]*kernel[3]+tmp[7424]*kernel[4]+tmp[7425]*kernel[5]+tmp[7523]*kernel[6]+tmp[7524]*kernel[7]+tmp[7525]*kernel[8];
				ans[7425]<=tmp[7324]*kernel[0]+tmp[7325]*kernel[1]+tmp[7326]*kernel[2]+tmp[7424]*kernel[3]+tmp[7425]*kernel[4]+tmp[7426]*kernel[5]+tmp[7524]*kernel[6]+tmp[7525]*kernel[7]+tmp[7526]*kernel[8];
				ans[7426]<=tmp[7325]*kernel[0]+tmp[7326]*kernel[1]+tmp[7327]*kernel[2]+tmp[7425]*kernel[3]+tmp[7426]*kernel[4]+tmp[7427]*kernel[5]+tmp[7525]*kernel[6]+tmp[7526]*kernel[7]+tmp[7527]*kernel[8];
				ans[7427]<=tmp[7326]*kernel[0]+tmp[7327]*kernel[1]+tmp[7328]*kernel[2]+tmp[7426]*kernel[3]+tmp[7427]*kernel[4]+tmp[7428]*kernel[5]+tmp[7526]*kernel[6]+tmp[7527]*kernel[7]+tmp[7528]*kernel[8];
				ans[7428]<=tmp[7327]*kernel[0]+tmp[7328]*kernel[1]+tmp[7329]*kernel[2]+tmp[7427]*kernel[3]+tmp[7428]*kernel[4]+tmp[7429]*kernel[5]+tmp[7527]*kernel[6]+tmp[7528]*kernel[7]+tmp[7529]*kernel[8];
				ans[7429]<=tmp[7328]*kernel[0]+tmp[7329]*kernel[1]+tmp[7330]*kernel[2]+tmp[7428]*kernel[3]+tmp[7429]*kernel[4]+tmp[7430]*kernel[5]+tmp[7528]*kernel[6]+tmp[7529]*kernel[7]+tmp[7530]*kernel[8];
				ans[7430]<=tmp[7329]*kernel[0]+tmp[7330]*kernel[1]+tmp[7331]*kernel[2]+tmp[7429]*kernel[3]+tmp[7430]*kernel[4]+tmp[7431]*kernel[5]+tmp[7529]*kernel[6]+tmp[7530]*kernel[7]+tmp[7531]*kernel[8];
				ans[7431]<=tmp[7330]*kernel[0]+tmp[7331]*kernel[1]+tmp[7332]*kernel[2]+tmp[7430]*kernel[3]+tmp[7431]*kernel[4]+tmp[7432]*kernel[5]+tmp[7530]*kernel[6]+tmp[7531]*kernel[7]+tmp[7532]*kernel[8];
				ans[7432]<=tmp[7331]*kernel[0]+tmp[7332]*kernel[1]+tmp[7333]*kernel[2]+tmp[7431]*kernel[3]+tmp[7432]*kernel[4]+tmp[7433]*kernel[5]+tmp[7531]*kernel[6]+tmp[7532]*kernel[7]+tmp[7533]*kernel[8];
				ans[7433]<=tmp[7332]*kernel[0]+tmp[7333]*kernel[1]+tmp[7334]*kernel[2]+tmp[7432]*kernel[3]+tmp[7433]*kernel[4]+tmp[7434]*kernel[5]+tmp[7532]*kernel[6]+tmp[7533]*kernel[7]+tmp[7534]*kernel[8];
				ans[7434]<=tmp[7333]*kernel[0]+tmp[7334]*kernel[1]+tmp[7335]*kernel[2]+tmp[7433]*kernel[3]+tmp[7434]*kernel[4]+tmp[7435]*kernel[5]+tmp[7533]*kernel[6]+tmp[7534]*kernel[7]+tmp[7535]*kernel[8];
				ans[7435]<=tmp[7334]*kernel[0]+tmp[7335]*kernel[1]+tmp[7336]*kernel[2]+tmp[7434]*kernel[3]+tmp[7435]*kernel[4]+tmp[7436]*kernel[5]+tmp[7534]*kernel[6]+tmp[7535]*kernel[7]+tmp[7536]*kernel[8];
				ans[7436]<=tmp[7335]*kernel[0]+tmp[7336]*kernel[1]+tmp[7337]*kernel[2]+tmp[7435]*kernel[3]+tmp[7436]*kernel[4]+tmp[7437]*kernel[5]+tmp[7535]*kernel[6]+tmp[7536]*kernel[7]+tmp[7537]*kernel[8];
				ans[7437]<=tmp[7336]*kernel[0]+tmp[7337]*kernel[1]+tmp[7338]*kernel[2]+tmp[7436]*kernel[3]+tmp[7437]*kernel[4]+tmp[7438]*kernel[5]+tmp[7536]*kernel[6]+tmp[7537]*kernel[7]+tmp[7538]*kernel[8];
				ans[7438]<=tmp[7337]*kernel[0]+tmp[7338]*kernel[1]+tmp[7339]*kernel[2]+tmp[7437]*kernel[3]+tmp[7438]*kernel[4]+tmp[7439]*kernel[5]+tmp[7537]*kernel[6]+tmp[7538]*kernel[7]+tmp[7539]*kernel[8];
				ans[7439]<=tmp[7338]*kernel[0]+tmp[7339]*kernel[1]+tmp[7340]*kernel[2]+tmp[7438]*kernel[3]+tmp[7439]*kernel[4]+tmp[7440]*kernel[5]+tmp[7538]*kernel[6]+tmp[7539]*kernel[7]+tmp[7540]*kernel[8];
				ans[7440]<=tmp[7339]*kernel[0]+tmp[7340]*kernel[1]+tmp[7341]*kernel[2]+tmp[7439]*kernel[3]+tmp[7440]*kernel[4]+tmp[7441]*kernel[5]+tmp[7539]*kernel[6]+tmp[7540]*kernel[7]+tmp[7541]*kernel[8];
				ans[7441]<=tmp[7340]*kernel[0]+tmp[7341]*kernel[1]+tmp[7342]*kernel[2]+tmp[7440]*kernel[3]+tmp[7441]*kernel[4]+tmp[7442]*kernel[5]+tmp[7540]*kernel[6]+tmp[7541]*kernel[7]+tmp[7542]*kernel[8];
				ans[7442]<=tmp[7341]*kernel[0]+tmp[7342]*kernel[1]+tmp[7343]*kernel[2]+tmp[7441]*kernel[3]+tmp[7442]*kernel[4]+tmp[7443]*kernel[5]+tmp[7541]*kernel[6]+tmp[7542]*kernel[7]+tmp[7543]*kernel[8];
				ans[7443]<=tmp[7342]*kernel[0]+tmp[7343]*kernel[1]+tmp[7344]*kernel[2]+tmp[7442]*kernel[3]+tmp[7443]*kernel[4]+tmp[7444]*kernel[5]+tmp[7542]*kernel[6]+tmp[7543]*kernel[7]+tmp[7544]*kernel[8];
				ans[7444]<=tmp[7343]*kernel[0]+tmp[7344]*kernel[1]+tmp[7345]*kernel[2]+tmp[7443]*kernel[3]+tmp[7444]*kernel[4]+tmp[7445]*kernel[5]+tmp[7543]*kernel[6]+tmp[7544]*kernel[7]+tmp[7545]*kernel[8];
				ans[7445]<=tmp[7344]*kernel[0]+tmp[7345]*kernel[1]+tmp[7346]*kernel[2]+tmp[7444]*kernel[3]+tmp[7445]*kernel[4]+tmp[7446]*kernel[5]+tmp[7544]*kernel[6]+tmp[7545]*kernel[7]+tmp[7546]*kernel[8];
				ans[7446]<=tmp[7345]*kernel[0]+tmp[7346]*kernel[1]+tmp[7347]*kernel[2]+tmp[7445]*kernel[3]+tmp[7446]*kernel[4]+tmp[7447]*kernel[5]+tmp[7545]*kernel[6]+tmp[7546]*kernel[7]+tmp[7547]*kernel[8];
				ans[7447]<=tmp[7346]*kernel[0]+tmp[7347]*kernel[1]+tmp[7348]*kernel[2]+tmp[7446]*kernel[3]+tmp[7447]*kernel[4]+tmp[7448]*kernel[5]+tmp[7546]*kernel[6]+tmp[7547]*kernel[7]+tmp[7548]*kernel[8];
				ans[7448]<=tmp[7347]*kernel[0]+tmp[7348]*kernel[1]+tmp[7349]*kernel[2]+tmp[7447]*kernel[3]+tmp[7448]*kernel[4]+tmp[7449]*kernel[5]+tmp[7547]*kernel[6]+tmp[7548]*kernel[7]+tmp[7549]*kernel[8];
				ans[7449]<=tmp[7348]*kernel[0]+tmp[7349]*kernel[1]+tmp[7350]*kernel[2]+tmp[7448]*kernel[3]+tmp[7449]*kernel[4]+tmp[7450]*kernel[5]+tmp[7548]*kernel[6]+tmp[7549]*kernel[7]+tmp[7550]*kernel[8];
				ans[7450]<=tmp[7349]*kernel[0]+tmp[7350]*kernel[1]+tmp[7351]*kernel[2]+tmp[7449]*kernel[3]+tmp[7450]*kernel[4]+tmp[7451]*kernel[5]+tmp[7549]*kernel[6]+tmp[7550]*kernel[7]+tmp[7551]*kernel[8];
				ans[7451]<=tmp[7350]*kernel[0]+tmp[7351]*kernel[1]+tmp[7352]*kernel[2]+tmp[7450]*kernel[3]+tmp[7451]*kernel[4]+tmp[7452]*kernel[5]+tmp[7550]*kernel[6]+tmp[7551]*kernel[7]+tmp[7552]*kernel[8];
				ans[7452]<=tmp[7351]*kernel[0]+tmp[7352]*kernel[1]+tmp[7353]*kernel[2]+tmp[7451]*kernel[3]+tmp[7452]*kernel[4]+tmp[7453]*kernel[5]+tmp[7551]*kernel[6]+tmp[7552]*kernel[7]+tmp[7553]*kernel[8];
				ans[7453]<=tmp[7352]*kernel[0]+tmp[7353]*kernel[1]+tmp[7354]*kernel[2]+tmp[7452]*kernel[3]+tmp[7453]*kernel[4]+tmp[7454]*kernel[5]+tmp[7552]*kernel[6]+tmp[7553]*kernel[7]+tmp[7554]*kernel[8];
				ans[7454]<=tmp[7353]*kernel[0]+tmp[7354]*kernel[1]+tmp[7355]*kernel[2]+tmp[7453]*kernel[3]+tmp[7454]*kernel[4]+tmp[7455]*kernel[5]+tmp[7553]*kernel[6]+tmp[7554]*kernel[7]+tmp[7555]*kernel[8];
				ans[7455]<=tmp[7354]*kernel[0]+tmp[7355]*kernel[1]+tmp[7356]*kernel[2]+tmp[7454]*kernel[3]+tmp[7455]*kernel[4]+tmp[7456]*kernel[5]+tmp[7554]*kernel[6]+tmp[7555]*kernel[7]+tmp[7556]*kernel[8];
				ans[7456]<=tmp[7355]*kernel[0]+tmp[7356]*kernel[1]+tmp[7357]*kernel[2]+tmp[7455]*kernel[3]+tmp[7456]*kernel[4]+tmp[7457]*kernel[5]+tmp[7555]*kernel[6]+tmp[7556]*kernel[7]+tmp[7557]*kernel[8];
				ans[7457]<=tmp[7356]*kernel[0]+tmp[7357]*kernel[1]+tmp[7358]*kernel[2]+tmp[7456]*kernel[3]+tmp[7457]*kernel[4]+tmp[7458]*kernel[5]+tmp[7556]*kernel[6]+tmp[7557]*kernel[7]+tmp[7558]*kernel[8];
				ans[7458]<=tmp[7357]*kernel[0]+tmp[7358]*kernel[1]+tmp[7359]*kernel[2]+tmp[7457]*kernel[3]+tmp[7458]*kernel[4]+tmp[7459]*kernel[5]+tmp[7557]*kernel[6]+tmp[7558]*kernel[7]+tmp[7559]*kernel[8];
				ans[7459]<=tmp[7358]*kernel[0]+tmp[7359]*kernel[1]+tmp[7360]*kernel[2]+tmp[7458]*kernel[3]+tmp[7459]*kernel[4]+tmp[7460]*kernel[5]+tmp[7558]*kernel[6]+tmp[7559]*kernel[7]+tmp[7560]*kernel[8];
				ans[7460]<=tmp[7359]*kernel[0]+tmp[7360]*kernel[1]+tmp[7361]*kernel[2]+tmp[7459]*kernel[3]+tmp[7460]*kernel[4]+tmp[7461]*kernel[5]+tmp[7559]*kernel[6]+tmp[7560]*kernel[7]+tmp[7561]*kernel[8];
				ans[7461]<=tmp[7360]*kernel[0]+tmp[7361]*kernel[1]+tmp[7362]*kernel[2]+tmp[7460]*kernel[3]+tmp[7461]*kernel[4]+tmp[7462]*kernel[5]+tmp[7560]*kernel[6]+tmp[7561]*kernel[7]+tmp[7562]*kernel[8];
				ans[7462]<=tmp[7361]*kernel[0]+tmp[7362]*kernel[1]+tmp[7363]*kernel[2]+tmp[7461]*kernel[3]+tmp[7462]*kernel[4]+tmp[7463]*kernel[5]+tmp[7561]*kernel[6]+tmp[7562]*kernel[7]+tmp[7563]*kernel[8];
				ans[7463]<=tmp[7362]*kernel[0]+tmp[7363]*kernel[1]+tmp[7364]*kernel[2]+tmp[7462]*kernel[3]+tmp[7463]*kernel[4]+tmp[7464]*kernel[5]+tmp[7562]*kernel[6]+tmp[7563]*kernel[7]+tmp[7564]*kernel[8];
				ans[7464]<=tmp[7363]*kernel[0]+tmp[7364]*kernel[1]+tmp[7365]*kernel[2]+tmp[7463]*kernel[3]+tmp[7464]*kernel[4]+tmp[7465]*kernel[5]+tmp[7563]*kernel[6]+tmp[7564]*kernel[7]+tmp[7565]*kernel[8];
				ans[7465]<=tmp[7364]*kernel[0]+tmp[7365]*kernel[1]+tmp[7366]*kernel[2]+tmp[7464]*kernel[3]+tmp[7465]*kernel[4]+tmp[7466]*kernel[5]+tmp[7564]*kernel[6]+tmp[7565]*kernel[7]+tmp[7566]*kernel[8];
				ans[7466]<=tmp[7365]*kernel[0]+tmp[7366]*kernel[1]+tmp[7367]*kernel[2]+tmp[7465]*kernel[3]+tmp[7466]*kernel[4]+tmp[7467]*kernel[5]+tmp[7565]*kernel[6]+tmp[7566]*kernel[7]+tmp[7567]*kernel[8];
				ans[7467]<=tmp[7366]*kernel[0]+tmp[7367]*kernel[1]+tmp[7368]*kernel[2]+tmp[7466]*kernel[3]+tmp[7467]*kernel[4]+tmp[7468]*kernel[5]+tmp[7566]*kernel[6]+tmp[7567]*kernel[7]+tmp[7568]*kernel[8];
				ans[7468]<=tmp[7367]*kernel[0]+tmp[7368]*kernel[1]+tmp[7369]*kernel[2]+tmp[7467]*kernel[3]+tmp[7468]*kernel[4]+tmp[7469]*kernel[5]+tmp[7567]*kernel[6]+tmp[7568]*kernel[7]+tmp[7569]*kernel[8];
				ans[7469]<=tmp[7368]*kernel[0]+tmp[7369]*kernel[1]+tmp[7370]*kernel[2]+tmp[7468]*kernel[3]+tmp[7469]*kernel[4]+tmp[7470]*kernel[5]+tmp[7568]*kernel[6]+tmp[7569]*kernel[7]+tmp[7570]*kernel[8];
				ans[7470]<=tmp[7369]*kernel[0]+tmp[7370]*kernel[1]+tmp[7371]*kernel[2]+tmp[7469]*kernel[3]+tmp[7470]*kernel[4]+tmp[7471]*kernel[5]+tmp[7569]*kernel[6]+tmp[7570]*kernel[7]+tmp[7571]*kernel[8];
				ans[7471]<=tmp[7370]*kernel[0]+tmp[7371]*kernel[1]+tmp[7372]*kernel[2]+tmp[7470]*kernel[3]+tmp[7471]*kernel[4]+tmp[7472]*kernel[5]+tmp[7570]*kernel[6]+tmp[7571]*kernel[7]+tmp[7572]*kernel[8];
				ans[7472]<=tmp[7371]*kernel[0]+tmp[7372]*kernel[1]+tmp[7373]*kernel[2]+tmp[7471]*kernel[3]+tmp[7472]*kernel[4]+tmp[7473]*kernel[5]+tmp[7571]*kernel[6]+tmp[7572]*kernel[7]+tmp[7573]*kernel[8];
				ans[7473]<=tmp[7372]*kernel[0]+tmp[7373]*kernel[1]+tmp[7374]*kernel[2]+tmp[7472]*kernel[3]+tmp[7473]*kernel[4]+tmp[7474]*kernel[5]+tmp[7572]*kernel[6]+tmp[7573]*kernel[7]+tmp[7574]*kernel[8];
				ans[7474]<=tmp[7373]*kernel[0]+tmp[7374]*kernel[1]+tmp[7375]*kernel[2]+tmp[7473]*kernel[3]+tmp[7474]*kernel[4]+tmp[7475]*kernel[5]+tmp[7573]*kernel[6]+tmp[7574]*kernel[7]+tmp[7575]*kernel[8];
				ans[7475]<=tmp[7374]*kernel[0]+tmp[7375]*kernel[1]+tmp[7376]*kernel[2]+tmp[7474]*kernel[3]+tmp[7475]*kernel[4]+tmp[7476]*kernel[5]+tmp[7574]*kernel[6]+tmp[7575]*kernel[7]+tmp[7576]*kernel[8];
				ans[7476]<=tmp[7375]*kernel[0]+tmp[7376]*kernel[1]+tmp[7377]*kernel[2]+tmp[7475]*kernel[3]+tmp[7476]*kernel[4]+tmp[7477]*kernel[5]+tmp[7575]*kernel[6]+tmp[7576]*kernel[7]+tmp[7577]*kernel[8];
				ans[7477]<=tmp[7376]*kernel[0]+tmp[7377]*kernel[1]+tmp[7378]*kernel[2]+tmp[7476]*kernel[3]+tmp[7477]*kernel[4]+tmp[7478]*kernel[5]+tmp[7576]*kernel[6]+tmp[7577]*kernel[7]+tmp[7578]*kernel[8];
				ans[7478]<=tmp[7377]*kernel[0]+tmp[7378]*kernel[1]+tmp[7379]*kernel[2]+tmp[7477]*kernel[3]+tmp[7478]*kernel[4]+tmp[7479]*kernel[5]+tmp[7577]*kernel[6]+tmp[7578]*kernel[7]+tmp[7579]*kernel[8];
				ans[7479]<=tmp[7378]*kernel[0]+tmp[7379]*kernel[1]+tmp[7380]*kernel[2]+tmp[7478]*kernel[3]+tmp[7479]*kernel[4]+tmp[7480]*kernel[5]+tmp[7578]*kernel[6]+tmp[7579]*kernel[7]+tmp[7580]*kernel[8];
				ans[7480]<=tmp[7379]*kernel[0]+tmp[7380]*kernel[1]+tmp[7381]*kernel[2]+tmp[7479]*kernel[3]+tmp[7480]*kernel[4]+tmp[7481]*kernel[5]+tmp[7579]*kernel[6]+tmp[7580]*kernel[7]+tmp[7581]*kernel[8];
				ans[7481]<=tmp[7380]*kernel[0]+tmp[7381]*kernel[1]+tmp[7382]*kernel[2]+tmp[7480]*kernel[3]+tmp[7481]*kernel[4]+tmp[7482]*kernel[5]+tmp[7580]*kernel[6]+tmp[7581]*kernel[7]+tmp[7582]*kernel[8];
				ans[7482]<=tmp[7381]*kernel[0]+tmp[7382]*kernel[1]+tmp[7383]*kernel[2]+tmp[7481]*kernel[3]+tmp[7482]*kernel[4]+tmp[7483]*kernel[5]+tmp[7581]*kernel[6]+tmp[7582]*kernel[7]+tmp[7583]*kernel[8];
				ans[7483]<=tmp[7382]*kernel[0]+tmp[7383]*kernel[1]+tmp[7384]*kernel[2]+tmp[7482]*kernel[3]+tmp[7483]*kernel[4]+tmp[7484]*kernel[5]+tmp[7582]*kernel[6]+tmp[7583]*kernel[7]+tmp[7584]*kernel[8];
				ans[7484]<=tmp[7383]*kernel[0]+tmp[7384]*kernel[1]+tmp[7385]*kernel[2]+tmp[7483]*kernel[3]+tmp[7484]*kernel[4]+tmp[7485]*kernel[5]+tmp[7583]*kernel[6]+tmp[7584]*kernel[7]+tmp[7585]*kernel[8];
				ans[7485]<=tmp[7384]*kernel[0]+tmp[7385]*kernel[1]+tmp[7386]*kernel[2]+tmp[7484]*kernel[3]+tmp[7485]*kernel[4]+tmp[7486]*kernel[5]+tmp[7584]*kernel[6]+tmp[7585]*kernel[7]+tmp[7586]*kernel[8];
				ans[7486]<=tmp[7385]*kernel[0]+tmp[7386]*kernel[1]+tmp[7387]*kernel[2]+tmp[7485]*kernel[3]+tmp[7486]*kernel[4]+tmp[7487]*kernel[5]+tmp[7585]*kernel[6]+tmp[7586]*kernel[7]+tmp[7587]*kernel[8];
				ans[7487]<=tmp[7386]*kernel[0]+tmp[7387]*kernel[1]+tmp[7388]*kernel[2]+tmp[7486]*kernel[3]+tmp[7487]*kernel[4]+tmp[7488]*kernel[5]+tmp[7586]*kernel[6]+tmp[7587]*kernel[7]+tmp[7588]*kernel[8];
				ans[7488]<=tmp[7387]*kernel[0]+tmp[7388]*kernel[1]+tmp[7389]*kernel[2]+tmp[7487]*kernel[3]+tmp[7488]*kernel[4]+tmp[7489]*kernel[5]+tmp[7587]*kernel[6]+tmp[7588]*kernel[7]+tmp[7589]*kernel[8];
				ans[7489]<=tmp[7388]*kernel[0]+tmp[7389]*kernel[1]+tmp[7390]*kernel[2]+tmp[7488]*kernel[3]+tmp[7489]*kernel[4]+tmp[7490]*kernel[5]+tmp[7588]*kernel[6]+tmp[7589]*kernel[7]+tmp[7590]*kernel[8];
				ans[7490]<=tmp[7389]*kernel[0]+tmp[7390]*kernel[1]+tmp[7391]*kernel[2]+tmp[7489]*kernel[3]+tmp[7490]*kernel[4]+tmp[7491]*kernel[5]+tmp[7589]*kernel[6]+tmp[7590]*kernel[7]+tmp[7591]*kernel[8];
				ans[7491]<=tmp[7390]*kernel[0]+tmp[7391]*kernel[1]+tmp[7392]*kernel[2]+tmp[7490]*kernel[3]+tmp[7491]*kernel[4]+tmp[7492]*kernel[5]+tmp[7590]*kernel[6]+tmp[7591]*kernel[7]+tmp[7592]*kernel[8];
				ans[7492]<=tmp[7391]*kernel[0]+tmp[7392]*kernel[1]+tmp[7393]*kernel[2]+tmp[7491]*kernel[3]+tmp[7492]*kernel[4]+tmp[7493]*kernel[5]+tmp[7591]*kernel[6]+tmp[7592]*kernel[7]+tmp[7593]*kernel[8];
				ans[7493]<=tmp[7392]*kernel[0]+tmp[7393]*kernel[1]+tmp[7394]*kernel[2]+tmp[7492]*kernel[3]+tmp[7493]*kernel[4]+tmp[7494]*kernel[5]+tmp[7592]*kernel[6]+tmp[7593]*kernel[7]+tmp[7594]*kernel[8];
				ans[7494]<=tmp[7393]*kernel[0]+tmp[7394]*kernel[1]+tmp[7395]*kernel[2]+tmp[7493]*kernel[3]+tmp[7494]*kernel[4]+tmp[7495]*kernel[5]+tmp[7593]*kernel[6]+tmp[7594]*kernel[7]+tmp[7595]*kernel[8];
				ans[7495]<=tmp[7394]*kernel[0]+tmp[7395]*kernel[1]+tmp[7396]*kernel[2]+tmp[7494]*kernel[3]+tmp[7495]*kernel[4]+tmp[7496]*kernel[5]+tmp[7594]*kernel[6]+tmp[7595]*kernel[7]+tmp[7596]*kernel[8];
				ans[7496]<=tmp[7395]*kernel[0]+tmp[7396]*kernel[1]+tmp[7397]*kernel[2]+tmp[7495]*kernel[3]+tmp[7496]*kernel[4]+tmp[7497]*kernel[5]+tmp[7595]*kernel[6]+tmp[7596]*kernel[7]+tmp[7597]*kernel[8];
				ans[7497]<=tmp[7396]*kernel[0]+tmp[7397]*kernel[1]+tmp[7398]*kernel[2]+tmp[7496]*kernel[3]+tmp[7497]*kernel[4]+tmp[7498]*kernel[5]+tmp[7596]*kernel[6]+tmp[7597]*kernel[7]+tmp[7598]*kernel[8];
				ans[7498]<=tmp[7397]*kernel[0]+tmp[7398]*kernel[1]+tmp[7399]*kernel[2]+tmp[7497]*kernel[3]+tmp[7498]*kernel[4]+tmp[7499]*kernel[5]+tmp[7597]*kernel[6]+tmp[7598]*kernel[7]+tmp[7599]*kernel[8];
				ans[7499]<=tmp[7398]*kernel[0]+tmp[7399]*kernel[1]+tmp[7498]*kernel[3]+tmp[7499]*kernel[4]+tmp[7598]*kernel[6]+tmp[7599]*kernel[7];
				ans[7500]<=tmp[7400]*kernel[1]+tmp[7401]*kernel[2]+tmp[7500]*kernel[4]+tmp[7501]*kernel[5]+tmp[7600]*kernel[7]+tmp[7601]*kernel[8];
				ans[7501]<=tmp[7400]*kernel[0]+tmp[7401]*kernel[1]+tmp[7402]*kernel[2]+tmp[7500]*kernel[3]+tmp[7501]*kernel[4]+tmp[7502]*kernel[5]+tmp[7600]*kernel[6]+tmp[7601]*kernel[7]+tmp[7602]*kernel[8];
				ans[7502]<=tmp[7401]*kernel[0]+tmp[7402]*kernel[1]+tmp[7403]*kernel[2]+tmp[7501]*kernel[3]+tmp[7502]*kernel[4]+tmp[7503]*kernel[5]+tmp[7601]*kernel[6]+tmp[7602]*kernel[7]+tmp[7603]*kernel[8];
				ans[7503]<=tmp[7402]*kernel[0]+tmp[7403]*kernel[1]+tmp[7404]*kernel[2]+tmp[7502]*kernel[3]+tmp[7503]*kernel[4]+tmp[7504]*kernel[5]+tmp[7602]*kernel[6]+tmp[7603]*kernel[7]+tmp[7604]*kernel[8];
				ans[7504]<=tmp[7403]*kernel[0]+tmp[7404]*kernel[1]+tmp[7405]*kernel[2]+tmp[7503]*kernel[3]+tmp[7504]*kernel[4]+tmp[7505]*kernel[5]+tmp[7603]*kernel[6]+tmp[7604]*kernel[7]+tmp[7605]*kernel[8];
				ans[7505]<=tmp[7404]*kernel[0]+tmp[7405]*kernel[1]+tmp[7406]*kernel[2]+tmp[7504]*kernel[3]+tmp[7505]*kernel[4]+tmp[7506]*kernel[5]+tmp[7604]*kernel[6]+tmp[7605]*kernel[7]+tmp[7606]*kernel[8];
				ans[7506]<=tmp[7405]*kernel[0]+tmp[7406]*kernel[1]+tmp[7407]*kernel[2]+tmp[7505]*kernel[3]+tmp[7506]*kernel[4]+tmp[7507]*kernel[5]+tmp[7605]*kernel[6]+tmp[7606]*kernel[7]+tmp[7607]*kernel[8];
				ans[7507]<=tmp[7406]*kernel[0]+tmp[7407]*kernel[1]+tmp[7408]*kernel[2]+tmp[7506]*kernel[3]+tmp[7507]*kernel[4]+tmp[7508]*kernel[5]+tmp[7606]*kernel[6]+tmp[7607]*kernel[7]+tmp[7608]*kernel[8];
				ans[7508]<=tmp[7407]*kernel[0]+tmp[7408]*kernel[1]+tmp[7409]*kernel[2]+tmp[7507]*kernel[3]+tmp[7508]*kernel[4]+tmp[7509]*kernel[5]+tmp[7607]*kernel[6]+tmp[7608]*kernel[7]+tmp[7609]*kernel[8];
				ans[7509]<=tmp[7408]*kernel[0]+tmp[7409]*kernel[1]+tmp[7410]*kernel[2]+tmp[7508]*kernel[3]+tmp[7509]*kernel[4]+tmp[7510]*kernel[5]+tmp[7608]*kernel[6]+tmp[7609]*kernel[7]+tmp[7610]*kernel[8];
				ans[7510]<=tmp[7409]*kernel[0]+tmp[7410]*kernel[1]+tmp[7411]*kernel[2]+tmp[7509]*kernel[3]+tmp[7510]*kernel[4]+tmp[7511]*kernel[5]+tmp[7609]*kernel[6]+tmp[7610]*kernel[7]+tmp[7611]*kernel[8];
				ans[7511]<=tmp[7410]*kernel[0]+tmp[7411]*kernel[1]+tmp[7412]*kernel[2]+tmp[7510]*kernel[3]+tmp[7511]*kernel[4]+tmp[7512]*kernel[5]+tmp[7610]*kernel[6]+tmp[7611]*kernel[7]+tmp[7612]*kernel[8];
				ans[7512]<=tmp[7411]*kernel[0]+tmp[7412]*kernel[1]+tmp[7413]*kernel[2]+tmp[7511]*kernel[3]+tmp[7512]*kernel[4]+tmp[7513]*kernel[5]+tmp[7611]*kernel[6]+tmp[7612]*kernel[7]+tmp[7613]*kernel[8];
				ans[7513]<=tmp[7412]*kernel[0]+tmp[7413]*kernel[1]+tmp[7414]*kernel[2]+tmp[7512]*kernel[3]+tmp[7513]*kernel[4]+tmp[7514]*kernel[5]+tmp[7612]*kernel[6]+tmp[7613]*kernel[7]+tmp[7614]*kernel[8];
				ans[7514]<=tmp[7413]*kernel[0]+tmp[7414]*kernel[1]+tmp[7415]*kernel[2]+tmp[7513]*kernel[3]+tmp[7514]*kernel[4]+tmp[7515]*kernel[5]+tmp[7613]*kernel[6]+tmp[7614]*kernel[7]+tmp[7615]*kernel[8];
				ans[7515]<=tmp[7414]*kernel[0]+tmp[7415]*kernel[1]+tmp[7416]*kernel[2]+tmp[7514]*kernel[3]+tmp[7515]*kernel[4]+tmp[7516]*kernel[5]+tmp[7614]*kernel[6]+tmp[7615]*kernel[7]+tmp[7616]*kernel[8];
				ans[7516]<=tmp[7415]*kernel[0]+tmp[7416]*kernel[1]+tmp[7417]*kernel[2]+tmp[7515]*kernel[3]+tmp[7516]*kernel[4]+tmp[7517]*kernel[5]+tmp[7615]*kernel[6]+tmp[7616]*kernel[7]+tmp[7617]*kernel[8];
				ans[7517]<=tmp[7416]*kernel[0]+tmp[7417]*kernel[1]+tmp[7418]*kernel[2]+tmp[7516]*kernel[3]+tmp[7517]*kernel[4]+tmp[7518]*kernel[5]+tmp[7616]*kernel[6]+tmp[7617]*kernel[7]+tmp[7618]*kernel[8];
				ans[7518]<=tmp[7417]*kernel[0]+tmp[7418]*kernel[1]+tmp[7419]*kernel[2]+tmp[7517]*kernel[3]+tmp[7518]*kernel[4]+tmp[7519]*kernel[5]+tmp[7617]*kernel[6]+tmp[7618]*kernel[7]+tmp[7619]*kernel[8];
				ans[7519]<=tmp[7418]*kernel[0]+tmp[7419]*kernel[1]+tmp[7420]*kernel[2]+tmp[7518]*kernel[3]+tmp[7519]*kernel[4]+tmp[7520]*kernel[5]+tmp[7618]*kernel[6]+tmp[7619]*kernel[7]+tmp[7620]*kernel[8];
				ans[7520]<=tmp[7419]*kernel[0]+tmp[7420]*kernel[1]+tmp[7421]*kernel[2]+tmp[7519]*kernel[3]+tmp[7520]*kernel[4]+tmp[7521]*kernel[5]+tmp[7619]*kernel[6]+tmp[7620]*kernel[7]+tmp[7621]*kernel[8];
				ans[7521]<=tmp[7420]*kernel[0]+tmp[7421]*kernel[1]+tmp[7422]*kernel[2]+tmp[7520]*kernel[3]+tmp[7521]*kernel[4]+tmp[7522]*kernel[5]+tmp[7620]*kernel[6]+tmp[7621]*kernel[7]+tmp[7622]*kernel[8];
				ans[7522]<=tmp[7421]*kernel[0]+tmp[7422]*kernel[1]+tmp[7423]*kernel[2]+tmp[7521]*kernel[3]+tmp[7522]*kernel[4]+tmp[7523]*kernel[5]+tmp[7621]*kernel[6]+tmp[7622]*kernel[7]+tmp[7623]*kernel[8];
				ans[7523]<=tmp[7422]*kernel[0]+tmp[7423]*kernel[1]+tmp[7424]*kernel[2]+tmp[7522]*kernel[3]+tmp[7523]*kernel[4]+tmp[7524]*kernel[5]+tmp[7622]*kernel[6]+tmp[7623]*kernel[7]+tmp[7624]*kernel[8];
				ans[7524]<=tmp[7423]*kernel[0]+tmp[7424]*kernel[1]+tmp[7425]*kernel[2]+tmp[7523]*kernel[3]+tmp[7524]*kernel[4]+tmp[7525]*kernel[5]+tmp[7623]*kernel[6]+tmp[7624]*kernel[7]+tmp[7625]*kernel[8];
				ans[7525]<=tmp[7424]*kernel[0]+tmp[7425]*kernel[1]+tmp[7426]*kernel[2]+tmp[7524]*kernel[3]+tmp[7525]*kernel[4]+tmp[7526]*kernel[5]+tmp[7624]*kernel[6]+tmp[7625]*kernel[7]+tmp[7626]*kernel[8];
				ans[7526]<=tmp[7425]*kernel[0]+tmp[7426]*kernel[1]+tmp[7427]*kernel[2]+tmp[7525]*kernel[3]+tmp[7526]*kernel[4]+tmp[7527]*kernel[5]+tmp[7625]*kernel[6]+tmp[7626]*kernel[7]+tmp[7627]*kernel[8];
				ans[7527]<=tmp[7426]*kernel[0]+tmp[7427]*kernel[1]+tmp[7428]*kernel[2]+tmp[7526]*kernel[3]+tmp[7527]*kernel[4]+tmp[7528]*kernel[5]+tmp[7626]*kernel[6]+tmp[7627]*kernel[7]+tmp[7628]*kernel[8];
				ans[7528]<=tmp[7427]*kernel[0]+tmp[7428]*kernel[1]+tmp[7429]*kernel[2]+tmp[7527]*kernel[3]+tmp[7528]*kernel[4]+tmp[7529]*kernel[5]+tmp[7627]*kernel[6]+tmp[7628]*kernel[7]+tmp[7629]*kernel[8];
				ans[7529]<=tmp[7428]*kernel[0]+tmp[7429]*kernel[1]+tmp[7430]*kernel[2]+tmp[7528]*kernel[3]+tmp[7529]*kernel[4]+tmp[7530]*kernel[5]+tmp[7628]*kernel[6]+tmp[7629]*kernel[7]+tmp[7630]*kernel[8];
				ans[7530]<=tmp[7429]*kernel[0]+tmp[7430]*kernel[1]+tmp[7431]*kernel[2]+tmp[7529]*kernel[3]+tmp[7530]*kernel[4]+tmp[7531]*kernel[5]+tmp[7629]*kernel[6]+tmp[7630]*kernel[7]+tmp[7631]*kernel[8];
				ans[7531]<=tmp[7430]*kernel[0]+tmp[7431]*kernel[1]+tmp[7432]*kernel[2]+tmp[7530]*kernel[3]+tmp[7531]*kernel[4]+tmp[7532]*kernel[5]+tmp[7630]*kernel[6]+tmp[7631]*kernel[7]+tmp[7632]*kernel[8];
				ans[7532]<=tmp[7431]*kernel[0]+tmp[7432]*kernel[1]+tmp[7433]*kernel[2]+tmp[7531]*kernel[3]+tmp[7532]*kernel[4]+tmp[7533]*kernel[5]+tmp[7631]*kernel[6]+tmp[7632]*kernel[7]+tmp[7633]*kernel[8];
				ans[7533]<=tmp[7432]*kernel[0]+tmp[7433]*kernel[1]+tmp[7434]*kernel[2]+tmp[7532]*kernel[3]+tmp[7533]*kernel[4]+tmp[7534]*kernel[5]+tmp[7632]*kernel[6]+tmp[7633]*kernel[7]+tmp[7634]*kernel[8];
				ans[7534]<=tmp[7433]*kernel[0]+tmp[7434]*kernel[1]+tmp[7435]*kernel[2]+tmp[7533]*kernel[3]+tmp[7534]*kernel[4]+tmp[7535]*kernel[5]+tmp[7633]*kernel[6]+tmp[7634]*kernel[7]+tmp[7635]*kernel[8];
				ans[7535]<=tmp[7434]*kernel[0]+tmp[7435]*kernel[1]+tmp[7436]*kernel[2]+tmp[7534]*kernel[3]+tmp[7535]*kernel[4]+tmp[7536]*kernel[5]+tmp[7634]*kernel[6]+tmp[7635]*kernel[7]+tmp[7636]*kernel[8];
				ans[7536]<=tmp[7435]*kernel[0]+tmp[7436]*kernel[1]+tmp[7437]*kernel[2]+tmp[7535]*kernel[3]+tmp[7536]*kernel[4]+tmp[7537]*kernel[5]+tmp[7635]*kernel[6]+tmp[7636]*kernel[7]+tmp[7637]*kernel[8];
				ans[7537]<=tmp[7436]*kernel[0]+tmp[7437]*kernel[1]+tmp[7438]*kernel[2]+tmp[7536]*kernel[3]+tmp[7537]*kernel[4]+tmp[7538]*kernel[5]+tmp[7636]*kernel[6]+tmp[7637]*kernel[7]+tmp[7638]*kernel[8];
				ans[7538]<=tmp[7437]*kernel[0]+tmp[7438]*kernel[1]+tmp[7439]*kernel[2]+tmp[7537]*kernel[3]+tmp[7538]*kernel[4]+tmp[7539]*kernel[5]+tmp[7637]*kernel[6]+tmp[7638]*kernel[7]+tmp[7639]*kernel[8];
				ans[7539]<=tmp[7438]*kernel[0]+tmp[7439]*kernel[1]+tmp[7440]*kernel[2]+tmp[7538]*kernel[3]+tmp[7539]*kernel[4]+tmp[7540]*kernel[5]+tmp[7638]*kernel[6]+tmp[7639]*kernel[7]+tmp[7640]*kernel[8];
				ans[7540]<=tmp[7439]*kernel[0]+tmp[7440]*kernel[1]+tmp[7441]*kernel[2]+tmp[7539]*kernel[3]+tmp[7540]*kernel[4]+tmp[7541]*kernel[5]+tmp[7639]*kernel[6]+tmp[7640]*kernel[7]+tmp[7641]*kernel[8];
				ans[7541]<=tmp[7440]*kernel[0]+tmp[7441]*kernel[1]+tmp[7442]*kernel[2]+tmp[7540]*kernel[3]+tmp[7541]*kernel[4]+tmp[7542]*kernel[5]+tmp[7640]*kernel[6]+tmp[7641]*kernel[7]+tmp[7642]*kernel[8];
				ans[7542]<=tmp[7441]*kernel[0]+tmp[7442]*kernel[1]+tmp[7443]*kernel[2]+tmp[7541]*kernel[3]+tmp[7542]*kernel[4]+tmp[7543]*kernel[5]+tmp[7641]*kernel[6]+tmp[7642]*kernel[7]+tmp[7643]*kernel[8];
				ans[7543]<=tmp[7442]*kernel[0]+tmp[7443]*kernel[1]+tmp[7444]*kernel[2]+tmp[7542]*kernel[3]+tmp[7543]*kernel[4]+tmp[7544]*kernel[5]+tmp[7642]*kernel[6]+tmp[7643]*kernel[7]+tmp[7644]*kernel[8];
				ans[7544]<=tmp[7443]*kernel[0]+tmp[7444]*kernel[1]+tmp[7445]*kernel[2]+tmp[7543]*kernel[3]+tmp[7544]*kernel[4]+tmp[7545]*kernel[5]+tmp[7643]*kernel[6]+tmp[7644]*kernel[7]+tmp[7645]*kernel[8];
				ans[7545]<=tmp[7444]*kernel[0]+tmp[7445]*kernel[1]+tmp[7446]*kernel[2]+tmp[7544]*kernel[3]+tmp[7545]*kernel[4]+tmp[7546]*kernel[5]+tmp[7644]*kernel[6]+tmp[7645]*kernel[7]+tmp[7646]*kernel[8];
				ans[7546]<=tmp[7445]*kernel[0]+tmp[7446]*kernel[1]+tmp[7447]*kernel[2]+tmp[7545]*kernel[3]+tmp[7546]*kernel[4]+tmp[7547]*kernel[5]+tmp[7645]*kernel[6]+tmp[7646]*kernel[7]+tmp[7647]*kernel[8];
				ans[7547]<=tmp[7446]*kernel[0]+tmp[7447]*kernel[1]+tmp[7448]*kernel[2]+tmp[7546]*kernel[3]+tmp[7547]*kernel[4]+tmp[7548]*kernel[5]+tmp[7646]*kernel[6]+tmp[7647]*kernel[7]+tmp[7648]*kernel[8];
				ans[7548]<=tmp[7447]*kernel[0]+tmp[7448]*kernel[1]+tmp[7449]*kernel[2]+tmp[7547]*kernel[3]+tmp[7548]*kernel[4]+tmp[7549]*kernel[5]+tmp[7647]*kernel[6]+tmp[7648]*kernel[7]+tmp[7649]*kernel[8];
				ans[7549]<=tmp[7448]*kernel[0]+tmp[7449]*kernel[1]+tmp[7450]*kernel[2]+tmp[7548]*kernel[3]+tmp[7549]*kernel[4]+tmp[7550]*kernel[5]+tmp[7648]*kernel[6]+tmp[7649]*kernel[7]+tmp[7650]*kernel[8];
				ans[7550]<=tmp[7449]*kernel[0]+tmp[7450]*kernel[1]+tmp[7451]*kernel[2]+tmp[7549]*kernel[3]+tmp[7550]*kernel[4]+tmp[7551]*kernel[5]+tmp[7649]*kernel[6]+tmp[7650]*kernel[7]+tmp[7651]*kernel[8];
				ans[7551]<=tmp[7450]*kernel[0]+tmp[7451]*kernel[1]+tmp[7452]*kernel[2]+tmp[7550]*kernel[3]+tmp[7551]*kernel[4]+tmp[7552]*kernel[5]+tmp[7650]*kernel[6]+tmp[7651]*kernel[7]+tmp[7652]*kernel[8];
				ans[7552]<=tmp[7451]*kernel[0]+tmp[7452]*kernel[1]+tmp[7453]*kernel[2]+tmp[7551]*kernel[3]+tmp[7552]*kernel[4]+tmp[7553]*kernel[5]+tmp[7651]*kernel[6]+tmp[7652]*kernel[7]+tmp[7653]*kernel[8];
				ans[7553]<=tmp[7452]*kernel[0]+tmp[7453]*kernel[1]+tmp[7454]*kernel[2]+tmp[7552]*kernel[3]+tmp[7553]*kernel[4]+tmp[7554]*kernel[5]+tmp[7652]*kernel[6]+tmp[7653]*kernel[7]+tmp[7654]*kernel[8];
				ans[7554]<=tmp[7453]*kernel[0]+tmp[7454]*kernel[1]+tmp[7455]*kernel[2]+tmp[7553]*kernel[3]+tmp[7554]*kernel[4]+tmp[7555]*kernel[5]+tmp[7653]*kernel[6]+tmp[7654]*kernel[7]+tmp[7655]*kernel[8];
				ans[7555]<=tmp[7454]*kernel[0]+tmp[7455]*kernel[1]+tmp[7456]*kernel[2]+tmp[7554]*kernel[3]+tmp[7555]*kernel[4]+tmp[7556]*kernel[5]+tmp[7654]*kernel[6]+tmp[7655]*kernel[7]+tmp[7656]*kernel[8];
				ans[7556]<=tmp[7455]*kernel[0]+tmp[7456]*kernel[1]+tmp[7457]*kernel[2]+tmp[7555]*kernel[3]+tmp[7556]*kernel[4]+tmp[7557]*kernel[5]+tmp[7655]*kernel[6]+tmp[7656]*kernel[7]+tmp[7657]*kernel[8];
				ans[7557]<=tmp[7456]*kernel[0]+tmp[7457]*kernel[1]+tmp[7458]*kernel[2]+tmp[7556]*kernel[3]+tmp[7557]*kernel[4]+tmp[7558]*kernel[5]+tmp[7656]*kernel[6]+tmp[7657]*kernel[7]+tmp[7658]*kernel[8];
				ans[7558]<=tmp[7457]*kernel[0]+tmp[7458]*kernel[1]+tmp[7459]*kernel[2]+tmp[7557]*kernel[3]+tmp[7558]*kernel[4]+tmp[7559]*kernel[5]+tmp[7657]*kernel[6]+tmp[7658]*kernel[7]+tmp[7659]*kernel[8];
				ans[7559]<=tmp[7458]*kernel[0]+tmp[7459]*kernel[1]+tmp[7460]*kernel[2]+tmp[7558]*kernel[3]+tmp[7559]*kernel[4]+tmp[7560]*kernel[5]+tmp[7658]*kernel[6]+tmp[7659]*kernel[7]+tmp[7660]*kernel[8];
				ans[7560]<=tmp[7459]*kernel[0]+tmp[7460]*kernel[1]+tmp[7461]*kernel[2]+tmp[7559]*kernel[3]+tmp[7560]*kernel[4]+tmp[7561]*kernel[5]+tmp[7659]*kernel[6]+tmp[7660]*kernel[7]+tmp[7661]*kernel[8];
				ans[7561]<=tmp[7460]*kernel[0]+tmp[7461]*kernel[1]+tmp[7462]*kernel[2]+tmp[7560]*kernel[3]+tmp[7561]*kernel[4]+tmp[7562]*kernel[5]+tmp[7660]*kernel[6]+tmp[7661]*kernel[7]+tmp[7662]*kernel[8];
				ans[7562]<=tmp[7461]*kernel[0]+tmp[7462]*kernel[1]+tmp[7463]*kernel[2]+tmp[7561]*kernel[3]+tmp[7562]*kernel[4]+tmp[7563]*kernel[5]+tmp[7661]*kernel[6]+tmp[7662]*kernel[7]+tmp[7663]*kernel[8];
				ans[7563]<=tmp[7462]*kernel[0]+tmp[7463]*kernel[1]+tmp[7464]*kernel[2]+tmp[7562]*kernel[3]+tmp[7563]*kernel[4]+tmp[7564]*kernel[5]+tmp[7662]*kernel[6]+tmp[7663]*kernel[7]+tmp[7664]*kernel[8];
				ans[7564]<=tmp[7463]*kernel[0]+tmp[7464]*kernel[1]+tmp[7465]*kernel[2]+tmp[7563]*kernel[3]+tmp[7564]*kernel[4]+tmp[7565]*kernel[5]+tmp[7663]*kernel[6]+tmp[7664]*kernel[7]+tmp[7665]*kernel[8];
				ans[7565]<=tmp[7464]*kernel[0]+tmp[7465]*kernel[1]+tmp[7466]*kernel[2]+tmp[7564]*kernel[3]+tmp[7565]*kernel[4]+tmp[7566]*kernel[5]+tmp[7664]*kernel[6]+tmp[7665]*kernel[7]+tmp[7666]*kernel[8];
				ans[7566]<=tmp[7465]*kernel[0]+tmp[7466]*kernel[1]+tmp[7467]*kernel[2]+tmp[7565]*kernel[3]+tmp[7566]*kernel[4]+tmp[7567]*kernel[5]+tmp[7665]*kernel[6]+tmp[7666]*kernel[7]+tmp[7667]*kernel[8];
				ans[7567]<=tmp[7466]*kernel[0]+tmp[7467]*kernel[1]+tmp[7468]*kernel[2]+tmp[7566]*kernel[3]+tmp[7567]*kernel[4]+tmp[7568]*kernel[5]+tmp[7666]*kernel[6]+tmp[7667]*kernel[7]+tmp[7668]*kernel[8];
				ans[7568]<=tmp[7467]*kernel[0]+tmp[7468]*kernel[1]+tmp[7469]*kernel[2]+tmp[7567]*kernel[3]+tmp[7568]*kernel[4]+tmp[7569]*kernel[5]+tmp[7667]*kernel[6]+tmp[7668]*kernel[7]+tmp[7669]*kernel[8];
				ans[7569]<=tmp[7468]*kernel[0]+tmp[7469]*kernel[1]+tmp[7470]*kernel[2]+tmp[7568]*kernel[3]+tmp[7569]*kernel[4]+tmp[7570]*kernel[5]+tmp[7668]*kernel[6]+tmp[7669]*kernel[7]+tmp[7670]*kernel[8];
				ans[7570]<=tmp[7469]*kernel[0]+tmp[7470]*kernel[1]+tmp[7471]*kernel[2]+tmp[7569]*kernel[3]+tmp[7570]*kernel[4]+tmp[7571]*kernel[5]+tmp[7669]*kernel[6]+tmp[7670]*kernel[7]+tmp[7671]*kernel[8];
				ans[7571]<=tmp[7470]*kernel[0]+tmp[7471]*kernel[1]+tmp[7472]*kernel[2]+tmp[7570]*kernel[3]+tmp[7571]*kernel[4]+tmp[7572]*kernel[5]+tmp[7670]*kernel[6]+tmp[7671]*kernel[7]+tmp[7672]*kernel[8];
				ans[7572]<=tmp[7471]*kernel[0]+tmp[7472]*kernel[1]+tmp[7473]*kernel[2]+tmp[7571]*kernel[3]+tmp[7572]*kernel[4]+tmp[7573]*kernel[5]+tmp[7671]*kernel[6]+tmp[7672]*kernel[7]+tmp[7673]*kernel[8];
				ans[7573]<=tmp[7472]*kernel[0]+tmp[7473]*kernel[1]+tmp[7474]*kernel[2]+tmp[7572]*kernel[3]+tmp[7573]*kernel[4]+tmp[7574]*kernel[5]+tmp[7672]*kernel[6]+tmp[7673]*kernel[7]+tmp[7674]*kernel[8];
				ans[7574]<=tmp[7473]*kernel[0]+tmp[7474]*kernel[1]+tmp[7475]*kernel[2]+tmp[7573]*kernel[3]+tmp[7574]*kernel[4]+tmp[7575]*kernel[5]+tmp[7673]*kernel[6]+tmp[7674]*kernel[7]+tmp[7675]*kernel[8];
				ans[7575]<=tmp[7474]*kernel[0]+tmp[7475]*kernel[1]+tmp[7476]*kernel[2]+tmp[7574]*kernel[3]+tmp[7575]*kernel[4]+tmp[7576]*kernel[5]+tmp[7674]*kernel[6]+tmp[7675]*kernel[7]+tmp[7676]*kernel[8];
				ans[7576]<=tmp[7475]*kernel[0]+tmp[7476]*kernel[1]+tmp[7477]*kernel[2]+tmp[7575]*kernel[3]+tmp[7576]*kernel[4]+tmp[7577]*kernel[5]+tmp[7675]*kernel[6]+tmp[7676]*kernel[7]+tmp[7677]*kernel[8];
				ans[7577]<=tmp[7476]*kernel[0]+tmp[7477]*kernel[1]+tmp[7478]*kernel[2]+tmp[7576]*kernel[3]+tmp[7577]*kernel[4]+tmp[7578]*kernel[5]+tmp[7676]*kernel[6]+tmp[7677]*kernel[7]+tmp[7678]*kernel[8];
				ans[7578]<=tmp[7477]*kernel[0]+tmp[7478]*kernel[1]+tmp[7479]*kernel[2]+tmp[7577]*kernel[3]+tmp[7578]*kernel[4]+tmp[7579]*kernel[5]+tmp[7677]*kernel[6]+tmp[7678]*kernel[7]+tmp[7679]*kernel[8];
				ans[7579]<=tmp[7478]*kernel[0]+tmp[7479]*kernel[1]+tmp[7480]*kernel[2]+tmp[7578]*kernel[3]+tmp[7579]*kernel[4]+tmp[7580]*kernel[5]+tmp[7678]*kernel[6]+tmp[7679]*kernel[7]+tmp[7680]*kernel[8];
				ans[7580]<=tmp[7479]*kernel[0]+tmp[7480]*kernel[1]+tmp[7481]*kernel[2]+tmp[7579]*kernel[3]+tmp[7580]*kernel[4]+tmp[7581]*kernel[5]+tmp[7679]*kernel[6]+tmp[7680]*kernel[7]+tmp[7681]*kernel[8];
				ans[7581]<=tmp[7480]*kernel[0]+tmp[7481]*kernel[1]+tmp[7482]*kernel[2]+tmp[7580]*kernel[3]+tmp[7581]*kernel[4]+tmp[7582]*kernel[5]+tmp[7680]*kernel[6]+tmp[7681]*kernel[7]+tmp[7682]*kernel[8];
				ans[7582]<=tmp[7481]*kernel[0]+tmp[7482]*kernel[1]+tmp[7483]*kernel[2]+tmp[7581]*kernel[3]+tmp[7582]*kernel[4]+tmp[7583]*kernel[5]+tmp[7681]*kernel[6]+tmp[7682]*kernel[7]+tmp[7683]*kernel[8];
				ans[7583]<=tmp[7482]*kernel[0]+tmp[7483]*kernel[1]+tmp[7484]*kernel[2]+tmp[7582]*kernel[3]+tmp[7583]*kernel[4]+tmp[7584]*kernel[5]+tmp[7682]*kernel[6]+tmp[7683]*kernel[7]+tmp[7684]*kernel[8];
				ans[7584]<=tmp[7483]*kernel[0]+tmp[7484]*kernel[1]+tmp[7485]*kernel[2]+tmp[7583]*kernel[3]+tmp[7584]*kernel[4]+tmp[7585]*kernel[5]+tmp[7683]*kernel[6]+tmp[7684]*kernel[7]+tmp[7685]*kernel[8];
				ans[7585]<=tmp[7484]*kernel[0]+tmp[7485]*kernel[1]+tmp[7486]*kernel[2]+tmp[7584]*kernel[3]+tmp[7585]*kernel[4]+tmp[7586]*kernel[5]+tmp[7684]*kernel[6]+tmp[7685]*kernel[7]+tmp[7686]*kernel[8];
				ans[7586]<=tmp[7485]*kernel[0]+tmp[7486]*kernel[1]+tmp[7487]*kernel[2]+tmp[7585]*kernel[3]+tmp[7586]*kernel[4]+tmp[7587]*kernel[5]+tmp[7685]*kernel[6]+tmp[7686]*kernel[7]+tmp[7687]*kernel[8];
				ans[7587]<=tmp[7486]*kernel[0]+tmp[7487]*kernel[1]+tmp[7488]*kernel[2]+tmp[7586]*kernel[3]+tmp[7587]*kernel[4]+tmp[7588]*kernel[5]+tmp[7686]*kernel[6]+tmp[7687]*kernel[7]+tmp[7688]*kernel[8];
				ans[7588]<=tmp[7487]*kernel[0]+tmp[7488]*kernel[1]+tmp[7489]*kernel[2]+tmp[7587]*kernel[3]+tmp[7588]*kernel[4]+tmp[7589]*kernel[5]+tmp[7687]*kernel[6]+tmp[7688]*kernel[7]+tmp[7689]*kernel[8];
				ans[7589]<=tmp[7488]*kernel[0]+tmp[7489]*kernel[1]+tmp[7490]*kernel[2]+tmp[7588]*kernel[3]+tmp[7589]*kernel[4]+tmp[7590]*kernel[5]+tmp[7688]*kernel[6]+tmp[7689]*kernel[7]+tmp[7690]*kernel[8];
				ans[7590]<=tmp[7489]*kernel[0]+tmp[7490]*kernel[1]+tmp[7491]*kernel[2]+tmp[7589]*kernel[3]+tmp[7590]*kernel[4]+tmp[7591]*kernel[5]+tmp[7689]*kernel[6]+tmp[7690]*kernel[7]+tmp[7691]*kernel[8];
				ans[7591]<=tmp[7490]*kernel[0]+tmp[7491]*kernel[1]+tmp[7492]*kernel[2]+tmp[7590]*kernel[3]+tmp[7591]*kernel[4]+tmp[7592]*kernel[5]+tmp[7690]*kernel[6]+tmp[7691]*kernel[7]+tmp[7692]*kernel[8];
				ans[7592]<=tmp[7491]*kernel[0]+tmp[7492]*kernel[1]+tmp[7493]*kernel[2]+tmp[7591]*kernel[3]+tmp[7592]*kernel[4]+tmp[7593]*kernel[5]+tmp[7691]*kernel[6]+tmp[7692]*kernel[7]+tmp[7693]*kernel[8];
				ans[7593]<=tmp[7492]*kernel[0]+tmp[7493]*kernel[1]+tmp[7494]*kernel[2]+tmp[7592]*kernel[3]+tmp[7593]*kernel[4]+tmp[7594]*kernel[5]+tmp[7692]*kernel[6]+tmp[7693]*kernel[7]+tmp[7694]*kernel[8];
				ans[7594]<=tmp[7493]*kernel[0]+tmp[7494]*kernel[1]+tmp[7495]*kernel[2]+tmp[7593]*kernel[3]+tmp[7594]*kernel[4]+tmp[7595]*kernel[5]+tmp[7693]*kernel[6]+tmp[7694]*kernel[7]+tmp[7695]*kernel[8];
				ans[7595]<=tmp[7494]*kernel[0]+tmp[7495]*kernel[1]+tmp[7496]*kernel[2]+tmp[7594]*kernel[3]+tmp[7595]*kernel[4]+tmp[7596]*kernel[5]+tmp[7694]*kernel[6]+tmp[7695]*kernel[7]+tmp[7696]*kernel[8];
				ans[7596]<=tmp[7495]*kernel[0]+tmp[7496]*kernel[1]+tmp[7497]*kernel[2]+tmp[7595]*kernel[3]+tmp[7596]*kernel[4]+tmp[7597]*kernel[5]+tmp[7695]*kernel[6]+tmp[7696]*kernel[7]+tmp[7697]*kernel[8];
				ans[7597]<=tmp[7496]*kernel[0]+tmp[7497]*kernel[1]+tmp[7498]*kernel[2]+tmp[7596]*kernel[3]+tmp[7597]*kernel[4]+tmp[7598]*kernel[5]+tmp[7696]*kernel[6]+tmp[7697]*kernel[7]+tmp[7698]*kernel[8];
				ans[7598]<=tmp[7497]*kernel[0]+tmp[7498]*kernel[1]+tmp[7499]*kernel[2]+tmp[7597]*kernel[3]+tmp[7598]*kernel[4]+tmp[7599]*kernel[5]+tmp[7697]*kernel[6]+tmp[7698]*kernel[7]+tmp[7699]*kernel[8];
				ans[7599]<=tmp[7498]*kernel[0]+tmp[7499]*kernel[1]+tmp[7598]*kernel[3]+tmp[7599]*kernel[4]+tmp[7698]*kernel[6]+tmp[7699]*kernel[7];
				ans[7600]<=tmp[7500]*kernel[1]+tmp[7501]*kernel[2]+tmp[7600]*kernel[4]+tmp[7601]*kernel[5]+tmp[7700]*kernel[7]+tmp[7701]*kernel[8];
				ans[7601]<=tmp[7500]*kernel[0]+tmp[7501]*kernel[1]+tmp[7502]*kernel[2]+tmp[7600]*kernel[3]+tmp[7601]*kernel[4]+tmp[7602]*kernel[5]+tmp[7700]*kernel[6]+tmp[7701]*kernel[7]+tmp[7702]*kernel[8];
				ans[7602]<=tmp[7501]*kernel[0]+tmp[7502]*kernel[1]+tmp[7503]*kernel[2]+tmp[7601]*kernel[3]+tmp[7602]*kernel[4]+tmp[7603]*kernel[5]+tmp[7701]*kernel[6]+tmp[7702]*kernel[7]+tmp[7703]*kernel[8];
				ans[7603]<=tmp[7502]*kernel[0]+tmp[7503]*kernel[1]+tmp[7504]*kernel[2]+tmp[7602]*kernel[3]+tmp[7603]*kernel[4]+tmp[7604]*kernel[5]+tmp[7702]*kernel[6]+tmp[7703]*kernel[7]+tmp[7704]*kernel[8];
				ans[7604]<=tmp[7503]*kernel[0]+tmp[7504]*kernel[1]+tmp[7505]*kernel[2]+tmp[7603]*kernel[3]+tmp[7604]*kernel[4]+tmp[7605]*kernel[5]+tmp[7703]*kernel[6]+tmp[7704]*kernel[7]+tmp[7705]*kernel[8];
				ans[7605]<=tmp[7504]*kernel[0]+tmp[7505]*kernel[1]+tmp[7506]*kernel[2]+tmp[7604]*kernel[3]+tmp[7605]*kernel[4]+tmp[7606]*kernel[5]+tmp[7704]*kernel[6]+tmp[7705]*kernel[7]+tmp[7706]*kernel[8];
				ans[7606]<=tmp[7505]*kernel[0]+tmp[7506]*kernel[1]+tmp[7507]*kernel[2]+tmp[7605]*kernel[3]+tmp[7606]*kernel[4]+tmp[7607]*kernel[5]+tmp[7705]*kernel[6]+tmp[7706]*kernel[7]+tmp[7707]*kernel[8];
				ans[7607]<=tmp[7506]*kernel[0]+tmp[7507]*kernel[1]+tmp[7508]*kernel[2]+tmp[7606]*kernel[3]+tmp[7607]*kernel[4]+tmp[7608]*kernel[5]+tmp[7706]*kernel[6]+tmp[7707]*kernel[7]+tmp[7708]*kernel[8];
				ans[7608]<=tmp[7507]*kernel[0]+tmp[7508]*kernel[1]+tmp[7509]*kernel[2]+tmp[7607]*kernel[3]+tmp[7608]*kernel[4]+tmp[7609]*kernel[5]+tmp[7707]*kernel[6]+tmp[7708]*kernel[7]+tmp[7709]*kernel[8];
				ans[7609]<=tmp[7508]*kernel[0]+tmp[7509]*kernel[1]+tmp[7510]*kernel[2]+tmp[7608]*kernel[3]+tmp[7609]*kernel[4]+tmp[7610]*kernel[5]+tmp[7708]*kernel[6]+tmp[7709]*kernel[7]+tmp[7710]*kernel[8];
				ans[7610]<=tmp[7509]*kernel[0]+tmp[7510]*kernel[1]+tmp[7511]*kernel[2]+tmp[7609]*kernel[3]+tmp[7610]*kernel[4]+tmp[7611]*kernel[5]+tmp[7709]*kernel[6]+tmp[7710]*kernel[7]+tmp[7711]*kernel[8];
				ans[7611]<=tmp[7510]*kernel[0]+tmp[7511]*kernel[1]+tmp[7512]*kernel[2]+tmp[7610]*kernel[3]+tmp[7611]*kernel[4]+tmp[7612]*kernel[5]+tmp[7710]*kernel[6]+tmp[7711]*kernel[7]+tmp[7712]*kernel[8];
				ans[7612]<=tmp[7511]*kernel[0]+tmp[7512]*kernel[1]+tmp[7513]*kernel[2]+tmp[7611]*kernel[3]+tmp[7612]*kernel[4]+tmp[7613]*kernel[5]+tmp[7711]*kernel[6]+tmp[7712]*kernel[7]+tmp[7713]*kernel[8];
				ans[7613]<=tmp[7512]*kernel[0]+tmp[7513]*kernel[1]+tmp[7514]*kernel[2]+tmp[7612]*kernel[3]+tmp[7613]*kernel[4]+tmp[7614]*kernel[5]+tmp[7712]*kernel[6]+tmp[7713]*kernel[7]+tmp[7714]*kernel[8];
				ans[7614]<=tmp[7513]*kernel[0]+tmp[7514]*kernel[1]+tmp[7515]*kernel[2]+tmp[7613]*kernel[3]+tmp[7614]*kernel[4]+tmp[7615]*kernel[5]+tmp[7713]*kernel[6]+tmp[7714]*kernel[7]+tmp[7715]*kernel[8];
				ans[7615]<=tmp[7514]*kernel[0]+tmp[7515]*kernel[1]+tmp[7516]*kernel[2]+tmp[7614]*kernel[3]+tmp[7615]*kernel[4]+tmp[7616]*kernel[5]+tmp[7714]*kernel[6]+tmp[7715]*kernel[7]+tmp[7716]*kernel[8];
				ans[7616]<=tmp[7515]*kernel[0]+tmp[7516]*kernel[1]+tmp[7517]*kernel[2]+tmp[7615]*kernel[3]+tmp[7616]*kernel[4]+tmp[7617]*kernel[5]+tmp[7715]*kernel[6]+tmp[7716]*kernel[7]+tmp[7717]*kernel[8];
				ans[7617]<=tmp[7516]*kernel[0]+tmp[7517]*kernel[1]+tmp[7518]*kernel[2]+tmp[7616]*kernel[3]+tmp[7617]*kernel[4]+tmp[7618]*kernel[5]+tmp[7716]*kernel[6]+tmp[7717]*kernel[7]+tmp[7718]*kernel[8];
				ans[7618]<=tmp[7517]*kernel[0]+tmp[7518]*kernel[1]+tmp[7519]*kernel[2]+tmp[7617]*kernel[3]+tmp[7618]*kernel[4]+tmp[7619]*kernel[5]+tmp[7717]*kernel[6]+tmp[7718]*kernel[7]+tmp[7719]*kernel[8];
				ans[7619]<=tmp[7518]*kernel[0]+tmp[7519]*kernel[1]+tmp[7520]*kernel[2]+tmp[7618]*kernel[3]+tmp[7619]*kernel[4]+tmp[7620]*kernel[5]+tmp[7718]*kernel[6]+tmp[7719]*kernel[7]+tmp[7720]*kernel[8];
				ans[7620]<=tmp[7519]*kernel[0]+tmp[7520]*kernel[1]+tmp[7521]*kernel[2]+tmp[7619]*kernel[3]+tmp[7620]*kernel[4]+tmp[7621]*kernel[5]+tmp[7719]*kernel[6]+tmp[7720]*kernel[7]+tmp[7721]*kernel[8];
				ans[7621]<=tmp[7520]*kernel[0]+tmp[7521]*kernel[1]+tmp[7522]*kernel[2]+tmp[7620]*kernel[3]+tmp[7621]*kernel[4]+tmp[7622]*kernel[5]+tmp[7720]*kernel[6]+tmp[7721]*kernel[7]+tmp[7722]*kernel[8];
				ans[7622]<=tmp[7521]*kernel[0]+tmp[7522]*kernel[1]+tmp[7523]*kernel[2]+tmp[7621]*kernel[3]+tmp[7622]*kernel[4]+tmp[7623]*kernel[5]+tmp[7721]*kernel[6]+tmp[7722]*kernel[7]+tmp[7723]*kernel[8];
				ans[7623]<=tmp[7522]*kernel[0]+tmp[7523]*kernel[1]+tmp[7524]*kernel[2]+tmp[7622]*kernel[3]+tmp[7623]*kernel[4]+tmp[7624]*kernel[5]+tmp[7722]*kernel[6]+tmp[7723]*kernel[7]+tmp[7724]*kernel[8];
				ans[7624]<=tmp[7523]*kernel[0]+tmp[7524]*kernel[1]+tmp[7525]*kernel[2]+tmp[7623]*kernel[3]+tmp[7624]*kernel[4]+tmp[7625]*kernel[5]+tmp[7723]*kernel[6]+tmp[7724]*kernel[7]+tmp[7725]*kernel[8];
				ans[7625]<=tmp[7524]*kernel[0]+tmp[7525]*kernel[1]+tmp[7526]*kernel[2]+tmp[7624]*kernel[3]+tmp[7625]*kernel[4]+tmp[7626]*kernel[5]+tmp[7724]*kernel[6]+tmp[7725]*kernel[7]+tmp[7726]*kernel[8];
				ans[7626]<=tmp[7525]*kernel[0]+tmp[7526]*kernel[1]+tmp[7527]*kernel[2]+tmp[7625]*kernel[3]+tmp[7626]*kernel[4]+tmp[7627]*kernel[5]+tmp[7725]*kernel[6]+tmp[7726]*kernel[7]+tmp[7727]*kernel[8];
				ans[7627]<=tmp[7526]*kernel[0]+tmp[7527]*kernel[1]+tmp[7528]*kernel[2]+tmp[7626]*kernel[3]+tmp[7627]*kernel[4]+tmp[7628]*kernel[5]+tmp[7726]*kernel[6]+tmp[7727]*kernel[7]+tmp[7728]*kernel[8];
				ans[7628]<=tmp[7527]*kernel[0]+tmp[7528]*kernel[1]+tmp[7529]*kernel[2]+tmp[7627]*kernel[3]+tmp[7628]*kernel[4]+tmp[7629]*kernel[5]+tmp[7727]*kernel[6]+tmp[7728]*kernel[7]+tmp[7729]*kernel[8];
				ans[7629]<=tmp[7528]*kernel[0]+tmp[7529]*kernel[1]+tmp[7530]*kernel[2]+tmp[7628]*kernel[3]+tmp[7629]*kernel[4]+tmp[7630]*kernel[5]+tmp[7728]*kernel[6]+tmp[7729]*kernel[7]+tmp[7730]*kernel[8];
				ans[7630]<=tmp[7529]*kernel[0]+tmp[7530]*kernel[1]+tmp[7531]*kernel[2]+tmp[7629]*kernel[3]+tmp[7630]*kernel[4]+tmp[7631]*kernel[5]+tmp[7729]*kernel[6]+tmp[7730]*kernel[7]+tmp[7731]*kernel[8];
				ans[7631]<=tmp[7530]*kernel[0]+tmp[7531]*kernel[1]+tmp[7532]*kernel[2]+tmp[7630]*kernel[3]+tmp[7631]*kernel[4]+tmp[7632]*kernel[5]+tmp[7730]*kernel[6]+tmp[7731]*kernel[7]+tmp[7732]*kernel[8];
				ans[7632]<=tmp[7531]*kernel[0]+tmp[7532]*kernel[1]+tmp[7533]*kernel[2]+tmp[7631]*kernel[3]+tmp[7632]*kernel[4]+tmp[7633]*kernel[5]+tmp[7731]*kernel[6]+tmp[7732]*kernel[7]+tmp[7733]*kernel[8];
				ans[7633]<=tmp[7532]*kernel[0]+tmp[7533]*kernel[1]+tmp[7534]*kernel[2]+tmp[7632]*kernel[3]+tmp[7633]*kernel[4]+tmp[7634]*kernel[5]+tmp[7732]*kernel[6]+tmp[7733]*kernel[7]+tmp[7734]*kernel[8];
				ans[7634]<=tmp[7533]*kernel[0]+tmp[7534]*kernel[1]+tmp[7535]*kernel[2]+tmp[7633]*kernel[3]+tmp[7634]*kernel[4]+tmp[7635]*kernel[5]+tmp[7733]*kernel[6]+tmp[7734]*kernel[7]+tmp[7735]*kernel[8];
				ans[7635]<=tmp[7534]*kernel[0]+tmp[7535]*kernel[1]+tmp[7536]*kernel[2]+tmp[7634]*kernel[3]+tmp[7635]*kernel[4]+tmp[7636]*kernel[5]+tmp[7734]*kernel[6]+tmp[7735]*kernel[7]+tmp[7736]*kernel[8];
				ans[7636]<=tmp[7535]*kernel[0]+tmp[7536]*kernel[1]+tmp[7537]*kernel[2]+tmp[7635]*kernel[3]+tmp[7636]*kernel[4]+tmp[7637]*kernel[5]+tmp[7735]*kernel[6]+tmp[7736]*kernel[7]+tmp[7737]*kernel[8];
				ans[7637]<=tmp[7536]*kernel[0]+tmp[7537]*kernel[1]+tmp[7538]*kernel[2]+tmp[7636]*kernel[3]+tmp[7637]*kernel[4]+tmp[7638]*kernel[5]+tmp[7736]*kernel[6]+tmp[7737]*kernel[7]+tmp[7738]*kernel[8];
				ans[7638]<=tmp[7537]*kernel[0]+tmp[7538]*kernel[1]+tmp[7539]*kernel[2]+tmp[7637]*kernel[3]+tmp[7638]*kernel[4]+tmp[7639]*kernel[5]+tmp[7737]*kernel[6]+tmp[7738]*kernel[7]+tmp[7739]*kernel[8];
				ans[7639]<=tmp[7538]*kernel[0]+tmp[7539]*kernel[1]+tmp[7540]*kernel[2]+tmp[7638]*kernel[3]+tmp[7639]*kernel[4]+tmp[7640]*kernel[5]+tmp[7738]*kernel[6]+tmp[7739]*kernel[7]+tmp[7740]*kernel[8];
				ans[7640]<=tmp[7539]*kernel[0]+tmp[7540]*kernel[1]+tmp[7541]*kernel[2]+tmp[7639]*kernel[3]+tmp[7640]*kernel[4]+tmp[7641]*kernel[5]+tmp[7739]*kernel[6]+tmp[7740]*kernel[7]+tmp[7741]*kernel[8];
				ans[7641]<=tmp[7540]*kernel[0]+tmp[7541]*kernel[1]+tmp[7542]*kernel[2]+tmp[7640]*kernel[3]+tmp[7641]*kernel[4]+tmp[7642]*kernel[5]+tmp[7740]*kernel[6]+tmp[7741]*kernel[7]+tmp[7742]*kernel[8];
				ans[7642]<=tmp[7541]*kernel[0]+tmp[7542]*kernel[1]+tmp[7543]*kernel[2]+tmp[7641]*kernel[3]+tmp[7642]*kernel[4]+tmp[7643]*kernel[5]+tmp[7741]*kernel[6]+tmp[7742]*kernel[7]+tmp[7743]*kernel[8];
				ans[7643]<=tmp[7542]*kernel[0]+tmp[7543]*kernel[1]+tmp[7544]*kernel[2]+tmp[7642]*kernel[3]+tmp[7643]*kernel[4]+tmp[7644]*kernel[5]+tmp[7742]*kernel[6]+tmp[7743]*kernel[7]+tmp[7744]*kernel[8];
				ans[7644]<=tmp[7543]*kernel[0]+tmp[7544]*kernel[1]+tmp[7545]*kernel[2]+tmp[7643]*kernel[3]+tmp[7644]*kernel[4]+tmp[7645]*kernel[5]+tmp[7743]*kernel[6]+tmp[7744]*kernel[7]+tmp[7745]*kernel[8];
				ans[7645]<=tmp[7544]*kernel[0]+tmp[7545]*kernel[1]+tmp[7546]*kernel[2]+tmp[7644]*kernel[3]+tmp[7645]*kernel[4]+tmp[7646]*kernel[5]+tmp[7744]*kernel[6]+tmp[7745]*kernel[7]+tmp[7746]*kernel[8];
				ans[7646]<=tmp[7545]*kernel[0]+tmp[7546]*kernel[1]+tmp[7547]*kernel[2]+tmp[7645]*kernel[3]+tmp[7646]*kernel[4]+tmp[7647]*kernel[5]+tmp[7745]*kernel[6]+tmp[7746]*kernel[7]+tmp[7747]*kernel[8];
				ans[7647]<=tmp[7546]*kernel[0]+tmp[7547]*kernel[1]+tmp[7548]*kernel[2]+tmp[7646]*kernel[3]+tmp[7647]*kernel[4]+tmp[7648]*kernel[5]+tmp[7746]*kernel[6]+tmp[7747]*kernel[7]+tmp[7748]*kernel[8];
				ans[7648]<=tmp[7547]*kernel[0]+tmp[7548]*kernel[1]+tmp[7549]*kernel[2]+tmp[7647]*kernel[3]+tmp[7648]*kernel[4]+tmp[7649]*kernel[5]+tmp[7747]*kernel[6]+tmp[7748]*kernel[7]+tmp[7749]*kernel[8];
				ans[7649]<=tmp[7548]*kernel[0]+tmp[7549]*kernel[1]+tmp[7550]*kernel[2]+tmp[7648]*kernel[3]+tmp[7649]*kernel[4]+tmp[7650]*kernel[5]+tmp[7748]*kernel[6]+tmp[7749]*kernel[7]+tmp[7750]*kernel[8];
				ans[7650]<=tmp[7549]*kernel[0]+tmp[7550]*kernel[1]+tmp[7551]*kernel[2]+tmp[7649]*kernel[3]+tmp[7650]*kernel[4]+tmp[7651]*kernel[5]+tmp[7749]*kernel[6]+tmp[7750]*kernel[7]+tmp[7751]*kernel[8];
				ans[7651]<=tmp[7550]*kernel[0]+tmp[7551]*kernel[1]+tmp[7552]*kernel[2]+tmp[7650]*kernel[3]+tmp[7651]*kernel[4]+tmp[7652]*kernel[5]+tmp[7750]*kernel[6]+tmp[7751]*kernel[7]+tmp[7752]*kernel[8];
				ans[7652]<=tmp[7551]*kernel[0]+tmp[7552]*kernel[1]+tmp[7553]*kernel[2]+tmp[7651]*kernel[3]+tmp[7652]*kernel[4]+tmp[7653]*kernel[5]+tmp[7751]*kernel[6]+tmp[7752]*kernel[7]+tmp[7753]*kernel[8];
				ans[7653]<=tmp[7552]*kernel[0]+tmp[7553]*kernel[1]+tmp[7554]*kernel[2]+tmp[7652]*kernel[3]+tmp[7653]*kernel[4]+tmp[7654]*kernel[5]+tmp[7752]*kernel[6]+tmp[7753]*kernel[7]+tmp[7754]*kernel[8];
				ans[7654]<=tmp[7553]*kernel[0]+tmp[7554]*kernel[1]+tmp[7555]*kernel[2]+tmp[7653]*kernel[3]+tmp[7654]*kernel[4]+tmp[7655]*kernel[5]+tmp[7753]*kernel[6]+tmp[7754]*kernel[7]+tmp[7755]*kernel[8];
				ans[7655]<=tmp[7554]*kernel[0]+tmp[7555]*kernel[1]+tmp[7556]*kernel[2]+tmp[7654]*kernel[3]+tmp[7655]*kernel[4]+tmp[7656]*kernel[5]+tmp[7754]*kernel[6]+tmp[7755]*kernel[7]+tmp[7756]*kernel[8];
				ans[7656]<=tmp[7555]*kernel[0]+tmp[7556]*kernel[1]+tmp[7557]*kernel[2]+tmp[7655]*kernel[3]+tmp[7656]*kernel[4]+tmp[7657]*kernel[5]+tmp[7755]*kernel[6]+tmp[7756]*kernel[7]+tmp[7757]*kernel[8];
				ans[7657]<=tmp[7556]*kernel[0]+tmp[7557]*kernel[1]+tmp[7558]*kernel[2]+tmp[7656]*kernel[3]+tmp[7657]*kernel[4]+tmp[7658]*kernel[5]+tmp[7756]*kernel[6]+tmp[7757]*kernel[7]+tmp[7758]*kernel[8];
				ans[7658]<=tmp[7557]*kernel[0]+tmp[7558]*kernel[1]+tmp[7559]*kernel[2]+tmp[7657]*kernel[3]+tmp[7658]*kernel[4]+tmp[7659]*kernel[5]+tmp[7757]*kernel[6]+tmp[7758]*kernel[7]+tmp[7759]*kernel[8];
				ans[7659]<=tmp[7558]*kernel[0]+tmp[7559]*kernel[1]+tmp[7560]*kernel[2]+tmp[7658]*kernel[3]+tmp[7659]*kernel[4]+tmp[7660]*kernel[5]+tmp[7758]*kernel[6]+tmp[7759]*kernel[7]+tmp[7760]*kernel[8];
				ans[7660]<=tmp[7559]*kernel[0]+tmp[7560]*kernel[1]+tmp[7561]*kernel[2]+tmp[7659]*kernel[3]+tmp[7660]*kernel[4]+tmp[7661]*kernel[5]+tmp[7759]*kernel[6]+tmp[7760]*kernel[7]+tmp[7761]*kernel[8];
				ans[7661]<=tmp[7560]*kernel[0]+tmp[7561]*kernel[1]+tmp[7562]*kernel[2]+tmp[7660]*kernel[3]+tmp[7661]*kernel[4]+tmp[7662]*kernel[5]+tmp[7760]*kernel[6]+tmp[7761]*kernel[7]+tmp[7762]*kernel[8];
				ans[7662]<=tmp[7561]*kernel[0]+tmp[7562]*kernel[1]+tmp[7563]*kernel[2]+tmp[7661]*kernel[3]+tmp[7662]*kernel[4]+tmp[7663]*kernel[5]+tmp[7761]*kernel[6]+tmp[7762]*kernel[7]+tmp[7763]*kernel[8];
				ans[7663]<=tmp[7562]*kernel[0]+tmp[7563]*kernel[1]+tmp[7564]*kernel[2]+tmp[7662]*kernel[3]+tmp[7663]*kernel[4]+tmp[7664]*kernel[5]+tmp[7762]*kernel[6]+tmp[7763]*kernel[7]+tmp[7764]*kernel[8];
				ans[7664]<=tmp[7563]*kernel[0]+tmp[7564]*kernel[1]+tmp[7565]*kernel[2]+tmp[7663]*kernel[3]+tmp[7664]*kernel[4]+tmp[7665]*kernel[5]+tmp[7763]*kernel[6]+tmp[7764]*kernel[7]+tmp[7765]*kernel[8];
				ans[7665]<=tmp[7564]*kernel[0]+tmp[7565]*kernel[1]+tmp[7566]*kernel[2]+tmp[7664]*kernel[3]+tmp[7665]*kernel[4]+tmp[7666]*kernel[5]+tmp[7764]*kernel[6]+tmp[7765]*kernel[7]+tmp[7766]*kernel[8];
				ans[7666]<=tmp[7565]*kernel[0]+tmp[7566]*kernel[1]+tmp[7567]*kernel[2]+tmp[7665]*kernel[3]+tmp[7666]*kernel[4]+tmp[7667]*kernel[5]+tmp[7765]*kernel[6]+tmp[7766]*kernel[7]+tmp[7767]*kernel[8];
				ans[7667]<=tmp[7566]*kernel[0]+tmp[7567]*kernel[1]+tmp[7568]*kernel[2]+tmp[7666]*kernel[3]+tmp[7667]*kernel[4]+tmp[7668]*kernel[5]+tmp[7766]*kernel[6]+tmp[7767]*kernel[7]+tmp[7768]*kernel[8];
				ans[7668]<=tmp[7567]*kernel[0]+tmp[7568]*kernel[1]+tmp[7569]*kernel[2]+tmp[7667]*kernel[3]+tmp[7668]*kernel[4]+tmp[7669]*kernel[5]+tmp[7767]*kernel[6]+tmp[7768]*kernel[7]+tmp[7769]*kernel[8];
				ans[7669]<=tmp[7568]*kernel[0]+tmp[7569]*kernel[1]+tmp[7570]*kernel[2]+tmp[7668]*kernel[3]+tmp[7669]*kernel[4]+tmp[7670]*kernel[5]+tmp[7768]*kernel[6]+tmp[7769]*kernel[7]+tmp[7770]*kernel[8];
				ans[7670]<=tmp[7569]*kernel[0]+tmp[7570]*kernel[1]+tmp[7571]*kernel[2]+tmp[7669]*kernel[3]+tmp[7670]*kernel[4]+tmp[7671]*kernel[5]+tmp[7769]*kernel[6]+tmp[7770]*kernel[7]+tmp[7771]*kernel[8];
				ans[7671]<=tmp[7570]*kernel[0]+tmp[7571]*kernel[1]+tmp[7572]*kernel[2]+tmp[7670]*kernel[3]+tmp[7671]*kernel[4]+tmp[7672]*kernel[5]+tmp[7770]*kernel[6]+tmp[7771]*kernel[7]+tmp[7772]*kernel[8];
				ans[7672]<=tmp[7571]*kernel[0]+tmp[7572]*kernel[1]+tmp[7573]*kernel[2]+tmp[7671]*kernel[3]+tmp[7672]*kernel[4]+tmp[7673]*kernel[5]+tmp[7771]*kernel[6]+tmp[7772]*kernel[7]+tmp[7773]*kernel[8];
				ans[7673]<=tmp[7572]*kernel[0]+tmp[7573]*kernel[1]+tmp[7574]*kernel[2]+tmp[7672]*kernel[3]+tmp[7673]*kernel[4]+tmp[7674]*kernel[5]+tmp[7772]*kernel[6]+tmp[7773]*kernel[7]+tmp[7774]*kernel[8];
				ans[7674]<=tmp[7573]*kernel[0]+tmp[7574]*kernel[1]+tmp[7575]*kernel[2]+tmp[7673]*kernel[3]+tmp[7674]*kernel[4]+tmp[7675]*kernel[5]+tmp[7773]*kernel[6]+tmp[7774]*kernel[7]+tmp[7775]*kernel[8];
				ans[7675]<=tmp[7574]*kernel[0]+tmp[7575]*kernel[1]+tmp[7576]*kernel[2]+tmp[7674]*kernel[3]+tmp[7675]*kernel[4]+tmp[7676]*kernel[5]+tmp[7774]*kernel[6]+tmp[7775]*kernel[7]+tmp[7776]*kernel[8];
				ans[7676]<=tmp[7575]*kernel[0]+tmp[7576]*kernel[1]+tmp[7577]*kernel[2]+tmp[7675]*kernel[3]+tmp[7676]*kernel[4]+tmp[7677]*kernel[5]+tmp[7775]*kernel[6]+tmp[7776]*kernel[7]+tmp[7777]*kernel[8];
				ans[7677]<=tmp[7576]*kernel[0]+tmp[7577]*kernel[1]+tmp[7578]*kernel[2]+tmp[7676]*kernel[3]+tmp[7677]*kernel[4]+tmp[7678]*kernel[5]+tmp[7776]*kernel[6]+tmp[7777]*kernel[7]+tmp[7778]*kernel[8];
				ans[7678]<=tmp[7577]*kernel[0]+tmp[7578]*kernel[1]+tmp[7579]*kernel[2]+tmp[7677]*kernel[3]+tmp[7678]*kernel[4]+tmp[7679]*kernel[5]+tmp[7777]*kernel[6]+tmp[7778]*kernel[7]+tmp[7779]*kernel[8];
				ans[7679]<=tmp[7578]*kernel[0]+tmp[7579]*kernel[1]+tmp[7580]*kernel[2]+tmp[7678]*kernel[3]+tmp[7679]*kernel[4]+tmp[7680]*kernel[5]+tmp[7778]*kernel[6]+tmp[7779]*kernel[7]+tmp[7780]*kernel[8];
				ans[7680]<=tmp[7579]*kernel[0]+tmp[7580]*kernel[1]+tmp[7581]*kernel[2]+tmp[7679]*kernel[3]+tmp[7680]*kernel[4]+tmp[7681]*kernel[5]+tmp[7779]*kernel[6]+tmp[7780]*kernel[7]+tmp[7781]*kernel[8];
				ans[7681]<=tmp[7580]*kernel[0]+tmp[7581]*kernel[1]+tmp[7582]*kernel[2]+tmp[7680]*kernel[3]+tmp[7681]*kernel[4]+tmp[7682]*kernel[5]+tmp[7780]*kernel[6]+tmp[7781]*kernel[7]+tmp[7782]*kernel[8];
				ans[7682]<=tmp[7581]*kernel[0]+tmp[7582]*kernel[1]+tmp[7583]*kernel[2]+tmp[7681]*kernel[3]+tmp[7682]*kernel[4]+tmp[7683]*kernel[5]+tmp[7781]*kernel[6]+tmp[7782]*kernel[7]+tmp[7783]*kernel[8];
				ans[7683]<=tmp[7582]*kernel[0]+tmp[7583]*kernel[1]+tmp[7584]*kernel[2]+tmp[7682]*kernel[3]+tmp[7683]*kernel[4]+tmp[7684]*kernel[5]+tmp[7782]*kernel[6]+tmp[7783]*kernel[7]+tmp[7784]*kernel[8];
				ans[7684]<=tmp[7583]*kernel[0]+tmp[7584]*kernel[1]+tmp[7585]*kernel[2]+tmp[7683]*kernel[3]+tmp[7684]*kernel[4]+tmp[7685]*kernel[5]+tmp[7783]*kernel[6]+tmp[7784]*kernel[7]+tmp[7785]*kernel[8];
				ans[7685]<=tmp[7584]*kernel[0]+tmp[7585]*kernel[1]+tmp[7586]*kernel[2]+tmp[7684]*kernel[3]+tmp[7685]*kernel[4]+tmp[7686]*kernel[5]+tmp[7784]*kernel[6]+tmp[7785]*kernel[7]+tmp[7786]*kernel[8];
				ans[7686]<=tmp[7585]*kernel[0]+tmp[7586]*kernel[1]+tmp[7587]*kernel[2]+tmp[7685]*kernel[3]+tmp[7686]*kernel[4]+tmp[7687]*kernel[5]+tmp[7785]*kernel[6]+tmp[7786]*kernel[7]+tmp[7787]*kernel[8];
				ans[7687]<=tmp[7586]*kernel[0]+tmp[7587]*kernel[1]+tmp[7588]*kernel[2]+tmp[7686]*kernel[3]+tmp[7687]*kernel[4]+tmp[7688]*kernel[5]+tmp[7786]*kernel[6]+tmp[7787]*kernel[7]+tmp[7788]*kernel[8];
				ans[7688]<=tmp[7587]*kernel[0]+tmp[7588]*kernel[1]+tmp[7589]*kernel[2]+tmp[7687]*kernel[3]+tmp[7688]*kernel[4]+tmp[7689]*kernel[5]+tmp[7787]*kernel[6]+tmp[7788]*kernel[7]+tmp[7789]*kernel[8];
				ans[7689]<=tmp[7588]*kernel[0]+tmp[7589]*kernel[1]+tmp[7590]*kernel[2]+tmp[7688]*kernel[3]+tmp[7689]*kernel[4]+tmp[7690]*kernel[5]+tmp[7788]*kernel[6]+tmp[7789]*kernel[7]+tmp[7790]*kernel[8];
				ans[7690]<=tmp[7589]*kernel[0]+tmp[7590]*kernel[1]+tmp[7591]*kernel[2]+tmp[7689]*kernel[3]+tmp[7690]*kernel[4]+tmp[7691]*kernel[5]+tmp[7789]*kernel[6]+tmp[7790]*kernel[7]+tmp[7791]*kernel[8];
				ans[7691]<=tmp[7590]*kernel[0]+tmp[7591]*kernel[1]+tmp[7592]*kernel[2]+tmp[7690]*kernel[3]+tmp[7691]*kernel[4]+tmp[7692]*kernel[5]+tmp[7790]*kernel[6]+tmp[7791]*kernel[7]+tmp[7792]*kernel[8];
				ans[7692]<=tmp[7591]*kernel[0]+tmp[7592]*kernel[1]+tmp[7593]*kernel[2]+tmp[7691]*kernel[3]+tmp[7692]*kernel[4]+tmp[7693]*kernel[5]+tmp[7791]*kernel[6]+tmp[7792]*kernel[7]+tmp[7793]*kernel[8];
				ans[7693]<=tmp[7592]*kernel[0]+tmp[7593]*kernel[1]+tmp[7594]*kernel[2]+tmp[7692]*kernel[3]+tmp[7693]*kernel[4]+tmp[7694]*kernel[5]+tmp[7792]*kernel[6]+tmp[7793]*kernel[7]+tmp[7794]*kernel[8];
				ans[7694]<=tmp[7593]*kernel[0]+tmp[7594]*kernel[1]+tmp[7595]*kernel[2]+tmp[7693]*kernel[3]+tmp[7694]*kernel[4]+tmp[7695]*kernel[5]+tmp[7793]*kernel[6]+tmp[7794]*kernel[7]+tmp[7795]*kernel[8];
				ans[7695]<=tmp[7594]*kernel[0]+tmp[7595]*kernel[1]+tmp[7596]*kernel[2]+tmp[7694]*kernel[3]+tmp[7695]*kernel[4]+tmp[7696]*kernel[5]+tmp[7794]*kernel[6]+tmp[7795]*kernel[7]+tmp[7796]*kernel[8];
				ans[7696]<=tmp[7595]*kernel[0]+tmp[7596]*kernel[1]+tmp[7597]*kernel[2]+tmp[7695]*kernel[3]+tmp[7696]*kernel[4]+tmp[7697]*kernel[5]+tmp[7795]*kernel[6]+tmp[7796]*kernel[7]+tmp[7797]*kernel[8];
				ans[7697]<=tmp[7596]*kernel[0]+tmp[7597]*kernel[1]+tmp[7598]*kernel[2]+tmp[7696]*kernel[3]+tmp[7697]*kernel[4]+tmp[7698]*kernel[5]+tmp[7796]*kernel[6]+tmp[7797]*kernel[7]+tmp[7798]*kernel[8];
				ans[7698]<=tmp[7597]*kernel[0]+tmp[7598]*kernel[1]+tmp[7599]*kernel[2]+tmp[7697]*kernel[3]+tmp[7698]*kernel[4]+tmp[7699]*kernel[5]+tmp[7797]*kernel[6]+tmp[7798]*kernel[7]+tmp[7799]*kernel[8];
				ans[7699]<=tmp[7598]*kernel[0]+tmp[7599]*kernel[1]+tmp[7698]*kernel[3]+tmp[7699]*kernel[4]+tmp[7798]*kernel[6]+tmp[7799]*kernel[7];
				ans[7700]<=tmp[7600]*kernel[1]+tmp[7601]*kernel[2]+tmp[7700]*kernel[4]+tmp[7701]*kernel[5]+tmp[7800]*kernel[7]+tmp[7801]*kernel[8];
				ans[7701]<=tmp[7600]*kernel[0]+tmp[7601]*kernel[1]+tmp[7602]*kernel[2]+tmp[7700]*kernel[3]+tmp[7701]*kernel[4]+tmp[7702]*kernel[5]+tmp[7800]*kernel[6]+tmp[7801]*kernel[7]+tmp[7802]*kernel[8];
				ans[7702]<=tmp[7601]*kernel[0]+tmp[7602]*kernel[1]+tmp[7603]*kernel[2]+tmp[7701]*kernel[3]+tmp[7702]*kernel[4]+tmp[7703]*kernel[5]+tmp[7801]*kernel[6]+tmp[7802]*kernel[7]+tmp[7803]*kernel[8];
				ans[7703]<=tmp[7602]*kernel[0]+tmp[7603]*kernel[1]+tmp[7604]*kernel[2]+tmp[7702]*kernel[3]+tmp[7703]*kernel[4]+tmp[7704]*kernel[5]+tmp[7802]*kernel[6]+tmp[7803]*kernel[7]+tmp[7804]*kernel[8];
				ans[7704]<=tmp[7603]*kernel[0]+tmp[7604]*kernel[1]+tmp[7605]*kernel[2]+tmp[7703]*kernel[3]+tmp[7704]*kernel[4]+tmp[7705]*kernel[5]+tmp[7803]*kernel[6]+tmp[7804]*kernel[7]+tmp[7805]*kernel[8];
				ans[7705]<=tmp[7604]*kernel[0]+tmp[7605]*kernel[1]+tmp[7606]*kernel[2]+tmp[7704]*kernel[3]+tmp[7705]*kernel[4]+tmp[7706]*kernel[5]+tmp[7804]*kernel[6]+tmp[7805]*kernel[7]+tmp[7806]*kernel[8];
				ans[7706]<=tmp[7605]*kernel[0]+tmp[7606]*kernel[1]+tmp[7607]*kernel[2]+tmp[7705]*kernel[3]+tmp[7706]*kernel[4]+tmp[7707]*kernel[5]+tmp[7805]*kernel[6]+tmp[7806]*kernel[7]+tmp[7807]*kernel[8];
				ans[7707]<=tmp[7606]*kernel[0]+tmp[7607]*kernel[1]+tmp[7608]*kernel[2]+tmp[7706]*kernel[3]+tmp[7707]*kernel[4]+tmp[7708]*kernel[5]+tmp[7806]*kernel[6]+tmp[7807]*kernel[7]+tmp[7808]*kernel[8];
				ans[7708]<=tmp[7607]*kernel[0]+tmp[7608]*kernel[1]+tmp[7609]*kernel[2]+tmp[7707]*kernel[3]+tmp[7708]*kernel[4]+tmp[7709]*kernel[5]+tmp[7807]*kernel[6]+tmp[7808]*kernel[7]+tmp[7809]*kernel[8];
				ans[7709]<=tmp[7608]*kernel[0]+tmp[7609]*kernel[1]+tmp[7610]*kernel[2]+tmp[7708]*kernel[3]+tmp[7709]*kernel[4]+tmp[7710]*kernel[5]+tmp[7808]*kernel[6]+tmp[7809]*kernel[7]+tmp[7810]*kernel[8];
				ans[7710]<=tmp[7609]*kernel[0]+tmp[7610]*kernel[1]+tmp[7611]*kernel[2]+tmp[7709]*kernel[3]+tmp[7710]*kernel[4]+tmp[7711]*kernel[5]+tmp[7809]*kernel[6]+tmp[7810]*kernel[7]+tmp[7811]*kernel[8];
				ans[7711]<=tmp[7610]*kernel[0]+tmp[7611]*kernel[1]+tmp[7612]*kernel[2]+tmp[7710]*kernel[3]+tmp[7711]*kernel[4]+tmp[7712]*kernel[5]+tmp[7810]*kernel[6]+tmp[7811]*kernel[7]+tmp[7812]*kernel[8];
				ans[7712]<=tmp[7611]*kernel[0]+tmp[7612]*kernel[1]+tmp[7613]*kernel[2]+tmp[7711]*kernel[3]+tmp[7712]*kernel[4]+tmp[7713]*kernel[5]+tmp[7811]*kernel[6]+tmp[7812]*kernel[7]+tmp[7813]*kernel[8];
				ans[7713]<=tmp[7612]*kernel[0]+tmp[7613]*kernel[1]+tmp[7614]*kernel[2]+tmp[7712]*kernel[3]+tmp[7713]*kernel[4]+tmp[7714]*kernel[5]+tmp[7812]*kernel[6]+tmp[7813]*kernel[7]+tmp[7814]*kernel[8];
				ans[7714]<=tmp[7613]*kernel[0]+tmp[7614]*kernel[1]+tmp[7615]*kernel[2]+tmp[7713]*kernel[3]+tmp[7714]*kernel[4]+tmp[7715]*kernel[5]+tmp[7813]*kernel[6]+tmp[7814]*kernel[7]+tmp[7815]*kernel[8];
				ans[7715]<=tmp[7614]*kernel[0]+tmp[7615]*kernel[1]+tmp[7616]*kernel[2]+tmp[7714]*kernel[3]+tmp[7715]*kernel[4]+tmp[7716]*kernel[5]+tmp[7814]*kernel[6]+tmp[7815]*kernel[7]+tmp[7816]*kernel[8];
				ans[7716]<=tmp[7615]*kernel[0]+tmp[7616]*kernel[1]+tmp[7617]*kernel[2]+tmp[7715]*kernel[3]+tmp[7716]*kernel[4]+tmp[7717]*kernel[5]+tmp[7815]*kernel[6]+tmp[7816]*kernel[7]+tmp[7817]*kernel[8];
				ans[7717]<=tmp[7616]*kernel[0]+tmp[7617]*kernel[1]+tmp[7618]*kernel[2]+tmp[7716]*kernel[3]+tmp[7717]*kernel[4]+tmp[7718]*kernel[5]+tmp[7816]*kernel[6]+tmp[7817]*kernel[7]+tmp[7818]*kernel[8];
				ans[7718]<=tmp[7617]*kernel[0]+tmp[7618]*kernel[1]+tmp[7619]*kernel[2]+tmp[7717]*kernel[3]+tmp[7718]*kernel[4]+tmp[7719]*kernel[5]+tmp[7817]*kernel[6]+tmp[7818]*kernel[7]+tmp[7819]*kernel[8];
				ans[7719]<=tmp[7618]*kernel[0]+tmp[7619]*kernel[1]+tmp[7620]*kernel[2]+tmp[7718]*kernel[3]+tmp[7719]*kernel[4]+tmp[7720]*kernel[5]+tmp[7818]*kernel[6]+tmp[7819]*kernel[7]+tmp[7820]*kernel[8];
				ans[7720]<=tmp[7619]*kernel[0]+tmp[7620]*kernel[1]+tmp[7621]*kernel[2]+tmp[7719]*kernel[3]+tmp[7720]*kernel[4]+tmp[7721]*kernel[5]+tmp[7819]*kernel[6]+tmp[7820]*kernel[7]+tmp[7821]*kernel[8];
				ans[7721]<=tmp[7620]*kernel[0]+tmp[7621]*kernel[1]+tmp[7622]*kernel[2]+tmp[7720]*kernel[3]+tmp[7721]*kernel[4]+tmp[7722]*kernel[5]+tmp[7820]*kernel[6]+tmp[7821]*kernel[7]+tmp[7822]*kernel[8];
				ans[7722]<=tmp[7621]*kernel[0]+tmp[7622]*kernel[1]+tmp[7623]*kernel[2]+tmp[7721]*kernel[3]+tmp[7722]*kernel[4]+tmp[7723]*kernel[5]+tmp[7821]*kernel[6]+tmp[7822]*kernel[7]+tmp[7823]*kernel[8];
				ans[7723]<=tmp[7622]*kernel[0]+tmp[7623]*kernel[1]+tmp[7624]*kernel[2]+tmp[7722]*kernel[3]+tmp[7723]*kernel[4]+tmp[7724]*kernel[5]+tmp[7822]*kernel[6]+tmp[7823]*kernel[7]+tmp[7824]*kernel[8];
				ans[7724]<=tmp[7623]*kernel[0]+tmp[7624]*kernel[1]+tmp[7625]*kernel[2]+tmp[7723]*kernel[3]+tmp[7724]*kernel[4]+tmp[7725]*kernel[5]+tmp[7823]*kernel[6]+tmp[7824]*kernel[7]+tmp[7825]*kernel[8];
				ans[7725]<=tmp[7624]*kernel[0]+tmp[7625]*kernel[1]+tmp[7626]*kernel[2]+tmp[7724]*kernel[3]+tmp[7725]*kernel[4]+tmp[7726]*kernel[5]+tmp[7824]*kernel[6]+tmp[7825]*kernel[7]+tmp[7826]*kernel[8];
				ans[7726]<=tmp[7625]*kernel[0]+tmp[7626]*kernel[1]+tmp[7627]*kernel[2]+tmp[7725]*kernel[3]+tmp[7726]*kernel[4]+tmp[7727]*kernel[5]+tmp[7825]*kernel[6]+tmp[7826]*kernel[7]+tmp[7827]*kernel[8];
				ans[7727]<=tmp[7626]*kernel[0]+tmp[7627]*kernel[1]+tmp[7628]*kernel[2]+tmp[7726]*kernel[3]+tmp[7727]*kernel[4]+tmp[7728]*kernel[5]+tmp[7826]*kernel[6]+tmp[7827]*kernel[7]+tmp[7828]*kernel[8];
				ans[7728]<=tmp[7627]*kernel[0]+tmp[7628]*kernel[1]+tmp[7629]*kernel[2]+tmp[7727]*kernel[3]+tmp[7728]*kernel[4]+tmp[7729]*kernel[5]+tmp[7827]*kernel[6]+tmp[7828]*kernel[7]+tmp[7829]*kernel[8];
				ans[7729]<=tmp[7628]*kernel[0]+tmp[7629]*kernel[1]+tmp[7630]*kernel[2]+tmp[7728]*kernel[3]+tmp[7729]*kernel[4]+tmp[7730]*kernel[5]+tmp[7828]*kernel[6]+tmp[7829]*kernel[7]+tmp[7830]*kernel[8];
				ans[7730]<=tmp[7629]*kernel[0]+tmp[7630]*kernel[1]+tmp[7631]*kernel[2]+tmp[7729]*kernel[3]+tmp[7730]*kernel[4]+tmp[7731]*kernel[5]+tmp[7829]*kernel[6]+tmp[7830]*kernel[7]+tmp[7831]*kernel[8];
				ans[7731]<=tmp[7630]*kernel[0]+tmp[7631]*kernel[1]+tmp[7632]*kernel[2]+tmp[7730]*kernel[3]+tmp[7731]*kernel[4]+tmp[7732]*kernel[5]+tmp[7830]*kernel[6]+tmp[7831]*kernel[7]+tmp[7832]*kernel[8];
				ans[7732]<=tmp[7631]*kernel[0]+tmp[7632]*kernel[1]+tmp[7633]*kernel[2]+tmp[7731]*kernel[3]+tmp[7732]*kernel[4]+tmp[7733]*kernel[5]+tmp[7831]*kernel[6]+tmp[7832]*kernel[7]+tmp[7833]*kernel[8];
				ans[7733]<=tmp[7632]*kernel[0]+tmp[7633]*kernel[1]+tmp[7634]*kernel[2]+tmp[7732]*kernel[3]+tmp[7733]*kernel[4]+tmp[7734]*kernel[5]+tmp[7832]*kernel[6]+tmp[7833]*kernel[7]+tmp[7834]*kernel[8];
				ans[7734]<=tmp[7633]*kernel[0]+tmp[7634]*kernel[1]+tmp[7635]*kernel[2]+tmp[7733]*kernel[3]+tmp[7734]*kernel[4]+tmp[7735]*kernel[5]+tmp[7833]*kernel[6]+tmp[7834]*kernel[7]+tmp[7835]*kernel[8];
				ans[7735]<=tmp[7634]*kernel[0]+tmp[7635]*kernel[1]+tmp[7636]*kernel[2]+tmp[7734]*kernel[3]+tmp[7735]*kernel[4]+tmp[7736]*kernel[5]+tmp[7834]*kernel[6]+tmp[7835]*kernel[7]+tmp[7836]*kernel[8];
				ans[7736]<=tmp[7635]*kernel[0]+tmp[7636]*kernel[1]+tmp[7637]*kernel[2]+tmp[7735]*kernel[3]+tmp[7736]*kernel[4]+tmp[7737]*kernel[5]+tmp[7835]*kernel[6]+tmp[7836]*kernel[7]+tmp[7837]*kernel[8];
				ans[7737]<=tmp[7636]*kernel[0]+tmp[7637]*kernel[1]+tmp[7638]*kernel[2]+tmp[7736]*kernel[3]+tmp[7737]*kernel[4]+tmp[7738]*kernel[5]+tmp[7836]*kernel[6]+tmp[7837]*kernel[7]+tmp[7838]*kernel[8];
				ans[7738]<=tmp[7637]*kernel[0]+tmp[7638]*kernel[1]+tmp[7639]*kernel[2]+tmp[7737]*kernel[3]+tmp[7738]*kernel[4]+tmp[7739]*kernel[5]+tmp[7837]*kernel[6]+tmp[7838]*kernel[7]+tmp[7839]*kernel[8];
				ans[7739]<=tmp[7638]*kernel[0]+tmp[7639]*kernel[1]+tmp[7640]*kernel[2]+tmp[7738]*kernel[3]+tmp[7739]*kernel[4]+tmp[7740]*kernel[5]+tmp[7838]*kernel[6]+tmp[7839]*kernel[7]+tmp[7840]*kernel[8];
				ans[7740]<=tmp[7639]*kernel[0]+tmp[7640]*kernel[1]+tmp[7641]*kernel[2]+tmp[7739]*kernel[3]+tmp[7740]*kernel[4]+tmp[7741]*kernel[5]+tmp[7839]*kernel[6]+tmp[7840]*kernel[7]+tmp[7841]*kernel[8];
				ans[7741]<=tmp[7640]*kernel[0]+tmp[7641]*kernel[1]+tmp[7642]*kernel[2]+tmp[7740]*kernel[3]+tmp[7741]*kernel[4]+tmp[7742]*kernel[5]+tmp[7840]*kernel[6]+tmp[7841]*kernel[7]+tmp[7842]*kernel[8];
				ans[7742]<=tmp[7641]*kernel[0]+tmp[7642]*kernel[1]+tmp[7643]*kernel[2]+tmp[7741]*kernel[3]+tmp[7742]*kernel[4]+tmp[7743]*kernel[5]+tmp[7841]*kernel[6]+tmp[7842]*kernel[7]+tmp[7843]*kernel[8];
				ans[7743]<=tmp[7642]*kernel[0]+tmp[7643]*kernel[1]+tmp[7644]*kernel[2]+tmp[7742]*kernel[3]+tmp[7743]*kernel[4]+tmp[7744]*kernel[5]+tmp[7842]*kernel[6]+tmp[7843]*kernel[7]+tmp[7844]*kernel[8];
				ans[7744]<=tmp[7643]*kernel[0]+tmp[7644]*kernel[1]+tmp[7645]*kernel[2]+tmp[7743]*kernel[3]+tmp[7744]*kernel[4]+tmp[7745]*kernel[5]+tmp[7843]*kernel[6]+tmp[7844]*kernel[7]+tmp[7845]*kernel[8];
				ans[7745]<=tmp[7644]*kernel[0]+tmp[7645]*kernel[1]+tmp[7646]*kernel[2]+tmp[7744]*kernel[3]+tmp[7745]*kernel[4]+tmp[7746]*kernel[5]+tmp[7844]*kernel[6]+tmp[7845]*kernel[7]+tmp[7846]*kernel[8];
				ans[7746]<=tmp[7645]*kernel[0]+tmp[7646]*kernel[1]+tmp[7647]*kernel[2]+tmp[7745]*kernel[3]+tmp[7746]*kernel[4]+tmp[7747]*kernel[5]+tmp[7845]*kernel[6]+tmp[7846]*kernel[7]+tmp[7847]*kernel[8];
				ans[7747]<=tmp[7646]*kernel[0]+tmp[7647]*kernel[1]+tmp[7648]*kernel[2]+tmp[7746]*kernel[3]+tmp[7747]*kernel[4]+tmp[7748]*kernel[5]+tmp[7846]*kernel[6]+tmp[7847]*kernel[7]+tmp[7848]*kernel[8];
				ans[7748]<=tmp[7647]*kernel[0]+tmp[7648]*kernel[1]+tmp[7649]*kernel[2]+tmp[7747]*kernel[3]+tmp[7748]*kernel[4]+tmp[7749]*kernel[5]+tmp[7847]*kernel[6]+tmp[7848]*kernel[7]+tmp[7849]*kernel[8];
				ans[7749]<=tmp[7648]*kernel[0]+tmp[7649]*kernel[1]+tmp[7650]*kernel[2]+tmp[7748]*kernel[3]+tmp[7749]*kernel[4]+tmp[7750]*kernel[5]+tmp[7848]*kernel[6]+tmp[7849]*kernel[7]+tmp[7850]*kernel[8];
				ans[7750]<=tmp[7649]*kernel[0]+tmp[7650]*kernel[1]+tmp[7651]*kernel[2]+tmp[7749]*kernel[3]+tmp[7750]*kernel[4]+tmp[7751]*kernel[5]+tmp[7849]*kernel[6]+tmp[7850]*kernel[7]+tmp[7851]*kernel[8];
				ans[7751]<=tmp[7650]*kernel[0]+tmp[7651]*kernel[1]+tmp[7652]*kernel[2]+tmp[7750]*kernel[3]+tmp[7751]*kernel[4]+tmp[7752]*kernel[5]+tmp[7850]*kernel[6]+tmp[7851]*kernel[7]+tmp[7852]*kernel[8];
				ans[7752]<=tmp[7651]*kernel[0]+tmp[7652]*kernel[1]+tmp[7653]*kernel[2]+tmp[7751]*kernel[3]+tmp[7752]*kernel[4]+tmp[7753]*kernel[5]+tmp[7851]*kernel[6]+tmp[7852]*kernel[7]+tmp[7853]*kernel[8];
				ans[7753]<=tmp[7652]*kernel[0]+tmp[7653]*kernel[1]+tmp[7654]*kernel[2]+tmp[7752]*kernel[3]+tmp[7753]*kernel[4]+tmp[7754]*kernel[5]+tmp[7852]*kernel[6]+tmp[7853]*kernel[7]+tmp[7854]*kernel[8];
				ans[7754]<=tmp[7653]*kernel[0]+tmp[7654]*kernel[1]+tmp[7655]*kernel[2]+tmp[7753]*kernel[3]+tmp[7754]*kernel[4]+tmp[7755]*kernel[5]+tmp[7853]*kernel[6]+tmp[7854]*kernel[7]+tmp[7855]*kernel[8];
				ans[7755]<=tmp[7654]*kernel[0]+tmp[7655]*kernel[1]+tmp[7656]*kernel[2]+tmp[7754]*kernel[3]+tmp[7755]*kernel[4]+tmp[7756]*kernel[5]+tmp[7854]*kernel[6]+tmp[7855]*kernel[7]+tmp[7856]*kernel[8];
				ans[7756]<=tmp[7655]*kernel[0]+tmp[7656]*kernel[1]+tmp[7657]*kernel[2]+tmp[7755]*kernel[3]+tmp[7756]*kernel[4]+tmp[7757]*kernel[5]+tmp[7855]*kernel[6]+tmp[7856]*kernel[7]+tmp[7857]*kernel[8];
				ans[7757]<=tmp[7656]*kernel[0]+tmp[7657]*kernel[1]+tmp[7658]*kernel[2]+tmp[7756]*kernel[3]+tmp[7757]*kernel[4]+tmp[7758]*kernel[5]+tmp[7856]*kernel[6]+tmp[7857]*kernel[7]+tmp[7858]*kernel[8];
				ans[7758]<=tmp[7657]*kernel[0]+tmp[7658]*kernel[1]+tmp[7659]*kernel[2]+tmp[7757]*kernel[3]+tmp[7758]*kernel[4]+tmp[7759]*kernel[5]+tmp[7857]*kernel[6]+tmp[7858]*kernel[7]+tmp[7859]*kernel[8];
				ans[7759]<=tmp[7658]*kernel[0]+tmp[7659]*kernel[1]+tmp[7660]*kernel[2]+tmp[7758]*kernel[3]+tmp[7759]*kernel[4]+tmp[7760]*kernel[5]+tmp[7858]*kernel[6]+tmp[7859]*kernel[7]+tmp[7860]*kernel[8];
				ans[7760]<=tmp[7659]*kernel[0]+tmp[7660]*kernel[1]+tmp[7661]*kernel[2]+tmp[7759]*kernel[3]+tmp[7760]*kernel[4]+tmp[7761]*kernel[5]+tmp[7859]*kernel[6]+tmp[7860]*kernel[7]+tmp[7861]*kernel[8];
				ans[7761]<=tmp[7660]*kernel[0]+tmp[7661]*kernel[1]+tmp[7662]*kernel[2]+tmp[7760]*kernel[3]+tmp[7761]*kernel[4]+tmp[7762]*kernel[5]+tmp[7860]*kernel[6]+tmp[7861]*kernel[7]+tmp[7862]*kernel[8];
				ans[7762]<=tmp[7661]*kernel[0]+tmp[7662]*kernel[1]+tmp[7663]*kernel[2]+tmp[7761]*kernel[3]+tmp[7762]*kernel[4]+tmp[7763]*kernel[5]+tmp[7861]*kernel[6]+tmp[7862]*kernel[7]+tmp[7863]*kernel[8];
				ans[7763]<=tmp[7662]*kernel[0]+tmp[7663]*kernel[1]+tmp[7664]*kernel[2]+tmp[7762]*kernel[3]+tmp[7763]*kernel[4]+tmp[7764]*kernel[5]+tmp[7862]*kernel[6]+tmp[7863]*kernel[7]+tmp[7864]*kernel[8];
				ans[7764]<=tmp[7663]*kernel[0]+tmp[7664]*kernel[1]+tmp[7665]*kernel[2]+tmp[7763]*kernel[3]+tmp[7764]*kernel[4]+tmp[7765]*kernel[5]+tmp[7863]*kernel[6]+tmp[7864]*kernel[7]+tmp[7865]*kernel[8];
				ans[7765]<=tmp[7664]*kernel[0]+tmp[7665]*kernel[1]+tmp[7666]*kernel[2]+tmp[7764]*kernel[3]+tmp[7765]*kernel[4]+tmp[7766]*kernel[5]+tmp[7864]*kernel[6]+tmp[7865]*kernel[7]+tmp[7866]*kernel[8];
				ans[7766]<=tmp[7665]*kernel[0]+tmp[7666]*kernel[1]+tmp[7667]*kernel[2]+tmp[7765]*kernel[3]+tmp[7766]*kernel[4]+tmp[7767]*kernel[5]+tmp[7865]*kernel[6]+tmp[7866]*kernel[7]+tmp[7867]*kernel[8];
				ans[7767]<=tmp[7666]*kernel[0]+tmp[7667]*kernel[1]+tmp[7668]*kernel[2]+tmp[7766]*kernel[3]+tmp[7767]*kernel[4]+tmp[7768]*kernel[5]+tmp[7866]*kernel[6]+tmp[7867]*kernel[7]+tmp[7868]*kernel[8];
				ans[7768]<=tmp[7667]*kernel[0]+tmp[7668]*kernel[1]+tmp[7669]*kernel[2]+tmp[7767]*kernel[3]+tmp[7768]*kernel[4]+tmp[7769]*kernel[5]+tmp[7867]*kernel[6]+tmp[7868]*kernel[7]+tmp[7869]*kernel[8];
				ans[7769]<=tmp[7668]*kernel[0]+tmp[7669]*kernel[1]+tmp[7670]*kernel[2]+tmp[7768]*kernel[3]+tmp[7769]*kernel[4]+tmp[7770]*kernel[5]+tmp[7868]*kernel[6]+tmp[7869]*kernel[7]+tmp[7870]*kernel[8];
				ans[7770]<=tmp[7669]*kernel[0]+tmp[7670]*kernel[1]+tmp[7671]*kernel[2]+tmp[7769]*kernel[3]+tmp[7770]*kernel[4]+tmp[7771]*kernel[5]+tmp[7869]*kernel[6]+tmp[7870]*kernel[7]+tmp[7871]*kernel[8];
				ans[7771]<=tmp[7670]*kernel[0]+tmp[7671]*kernel[1]+tmp[7672]*kernel[2]+tmp[7770]*kernel[3]+tmp[7771]*kernel[4]+tmp[7772]*kernel[5]+tmp[7870]*kernel[6]+tmp[7871]*kernel[7]+tmp[7872]*kernel[8];
				ans[7772]<=tmp[7671]*kernel[0]+tmp[7672]*kernel[1]+tmp[7673]*kernel[2]+tmp[7771]*kernel[3]+tmp[7772]*kernel[4]+tmp[7773]*kernel[5]+tmp[7871]*kernel[6]+tmp[7872]*kernel[7]+tmp[7873]*kernel[8];
				ans[7773]<=tmp[7672]*kernel[0]+tmp[7673]*kernel[1]+tmp[7674]*kernel[2]+tmp[7772]*kernel[3]+tmp[7773]*kernel[4]+tmp[7774]*kernel[5]+tmp[7872]*kernel[6]+tmp[7873]*kernel[7]+tmp[7874]*kernel[8];
				ans[7774]<=tmp[7673]*kernel[0]+tmp[7674]*kernel[1]+tmp[7675]*kernel[2]+tmp[7773]*kernel[3]+tmp[7774]*kernel[4]+tmp[7775]*kernel[5]+tmp[7873]*kernel[6]+tmp[7874]*kernel[7]+tmp[7875]*kernel[8];
				ans[7775]<=tmp[7674]*kernel[0]+tmp[7675]*kernel[1]+tmp[7676]*kernel[2]+tmp[7774]*kernel[3]+tmp[7775]*kernel[4]+tmp[7776]*kernel[5]+tmp[7874]*kernel[6]+tmp[7875]*kernel[7]+tmp[7876]*kernel[8];
				ans[7776]<=tmp[7675]*kernel[0]+tmp[7676]*kernel[1]+tmp[7677]*kernel[2]+tmp[7775]*kernel[3]+tmp[7776]*kernel[4]+tmp[7777]*kernel[5]+tmp[7875]*kernel[6]+tmp[7876]*kernel[7]+tmp[7877]*kernel[8];
				ans[7777]<=tmp[7676]*kernel[0]+tmp[7677]*kernel[1]+tmp[7678]*kernel[2]+tmp[7776]*kernel[3]+tmp[7777]*kernel[4]+tmp[7778]*kernel[5]+tmp[7876]*kernel[6]+tmp[7877]*kernel[7]+tmp[7878]*kernel[8];
				ans[7778]<=tmp[7677]*kernel[0]+tmp[7678]*kernel[1]+tmp[7679]*kernel[2]+tmp[7777]*kernel[3]+tmp[7778]*kernel[4]+tmp[7779]*kernel[5]+tmp[7877]*kernel[6]+tmp[7878]*kernel[7]+tmp[7879]*kernel[8];
				ans[7779]<=tmp[7678]*kernel[0]+tmp[7679]*kernel[1]+tmp[7680]*kernel[2]+tmp[7778]*kernel[3]+tmp[7779]*kernel[4]+tmp[7780]*kernel[5]+tmp[7878]*kernel[6]+tmp[7879]*kernel[7]+tmp[7880]*kernel[8];
				ans[7780]<=tmp[7679]*kernel[0]+tmp[7680]*kernel[1]+tmp[7681]*kernel[2]+tmp[7779]*kernel[3]+tmp[7780]*kernel[4]+tmp[7781]*kernel[5]+tmp[7879]*kernel[6]+tmp[7880]*kernel[7]+tmp[7881]*kernel[8];
				ans[7781]<=tmp[7680]*kernel[0]+tmp[7681]*kernel[1]+tmp[7682]*kernel[2]+tmp[7780]*kernel[3]+tmp[7781]*kernel[4]+tmp[7782]*kernel[5]+tmp[7880]*kernel[6]+tmp[7881]*kernel[7]+tmp[7882]*kernel[8];
				ans[7782]<=tmp[7681]*kernel[0]+tmp[7682]*kernel[1]+tmp[7683]*kernel[2]+tmp[7781]*kernel[3]+tmp[7782]*kernel[4]+tmp[7783]*kernel[5]+tmp[7881]*kernel[6]+tmp[7882]*kernel[7]+tmp[7883]*kernel[8];
				ans[7783]<=tmp[7682]*kernel[0]+tmp[7683]*kernel[1]+tmp[7684]*kernel[2]+tmp[7782]*kernel[3]+tmp[7783]*kernel[4]+tmp[7784]*kernel[5]+tmp[7882]*kernel[6]+tmp[7883]*kernel[7]+tmp[7884]*kernel[8];
				ans[7784]<=tmp[7683]*kernel[0]+tmp[7684]*kernel[1]+tmp[7685]*kernel[2]+tmp[7783]*kernel[3]+tmp[7784]*kernel[4]+tmp[7785]*kernel[5]+tmp[7883]*kernel[6]+tmp[7884]*kernel[7]+tmp[7885]*kernel[8];
				ans[7785]<=tmp[7684]*kernel[0]+tmp[7685]*kernel[1]+tmp[7686]*kernel[2]+tmp[7784]*kernel[3]+tmp[7785]*kernel[4]+tmp[7786]*kernel[5]+tmp[7884]*kernel[6]+tmp[7885]*kernel[7]+tmp[7886]*kernel[8];
				ans[7786]<=tmp[7685]*kernel[0]+tmp[7686]*kernel[1]+tmp[7687]*kernel[2]+tmp[7785]*kernel[3]+tmp[7786]*kernel[4]+tmp[7787]*kernel[5]+tmp[7885]*kernel[6]+tmp[7886]*kernel[7]+tmp[7887]*kernel[8];
				ans[7787]<=tmp[7686]*kernel[0]+tmp[7687]*kernel[1]+tmp[7688]*kernel[2]+tmp[7786]*kernel[3]+tmp[7787]*kernel[4]+tmp[7788]*kernel[5]+tmp[7886]*kernel[6]+tmp[7887]*kernel[7]+tmp[7888]*kernel[8];
				ans[7788]<=tmp[7687]*kernel[0]+tmp[7688]*kernel[1]+tmp[7689]*kernel[2]+tmp[7787]*kernel[3]+tmp[7788]*kernel[4]+tmp[7789]*kernel[5]+tmp[7887]*kernel[6]+tmp[7888]*kernel[7]+tmp[7889]*kernel[8];
				ans[7789]<=tmp[7688]*kernel[0]+tmp[7689]*kernel[1]+tmp[7690]*kernel[2]+tmp[7788]*kernel[3]+tmp[7789]*kernel[4]+tmp[7790]*kernel[5]+tmp[7888]*kernel[6]+tmp[7889]*kernel[7]+tmp[7890]*kernel[8];
				ans[7790]<=tmp[7689]*kernel[0]+tmp[7690]*kernel[1]+tmp[7691]*kernel[2]+tmp[7789]*kernel[3]+tmp[7790]*kernel[4]+tmp[7791]*kernel[5]+tmp[7889]*kernel[6]+tmp[7890]*kernel[7]+tmp[7891]*kernel[8];
				ans[7791]<=tmp[7690]*kernel[0]+tmp[7691]*kernel[1]+tmp[7692]*kernel[2]+tmp[7790]*kernel[3]+tmp[7791]*kernel[4]+tmp[7792]*kernel[5]+tmp[7890]*kernel[6]+tmp[7891]*kernel[7]+tmp[7892]*kernel[8];
				ans[7792]<=tmp[7691]*kernel[0]+tmp[7692]*kernel[1]+tmp[7693]*kernel[2]+tmp[7791]*kernel[3]+tmp[7792]*kernel[4]+tmp[7793]*kernel[5]+tmp[7891]*kernel[6]+tmp[7892]*kernel[7]+tmp[7893]*kernel[8];
				ans[7793]<=tmp[7692]*kernel[0]+tmp[7693]*kernel[1]+tmp[7694]*kernel[2]+tmp[7792]*kernel[3]+tmp[7793]*kernel[4]+tmp[7794]*kernel[5]+tmp[7892]*kernel[6]+tmp[7893]*kernel[7]+tmp[7894]*kernel[8];
				ans[7794]<=tmp[7693]*kernel[0]+tmp[7694]*kernel[1]+tmp[7695]*kernel[2]+tmp[7793]*kernel[3]+tmp[7794]*kernel[4]+tmp[7795]*kernel[5]+tmp[7893]*kernel[6]+tmp[7894]*kernel[7]+tmp[7895]*kernel[8];
				ans[7795]<=tmp[7694]*kernel[0]+tmp[7695]*kernel[1]+tmp[7696]*kernel[2]+tmp[7794]*kernel[3]+tmp[7795]*kernel[4]+tmp[7796]*kernel[5]+tmp[7894]*kernel[6]+tmp[7895]*kernel[7]+tmp[7896]*kernel[8];
				ans[7796]<=tmp[7695]*kernel[0]+tmp[7696]*kernel[1]+tmp[7697]*kernel[2]+tmp[7795]*kernel[3]+tmp[7796]*kernel[4]+tmp[7797]*kernel[5]+tmp[7895]*kernel[6]+tmp[7896]*kernel[7]+tmp[7897]*kernel[8];
				ans[7797]<=tmp[7696]*kernel[0]+tmp[7697]*kernel[1]+tmp[7698]*kernel[2]+tmp[7796]*kernel[3]+tmp[7797]*kernel[4]+tmp[7798]*kernel[5]+tmp[7896]*kernel[6]+tmp[7897]*kernel[7]+tmp[7898]*kernel[8];
				ans[7798]<=tmp[7697]*kernel[0]+tmp[7698]*kernel[1]+tmp[7699]*kernel[2]+tmp[7797]*kernel[3]+tmp[7798]*kernel[4]+tmp[7799]*kernel[5]+tmp[7897]*kernel[6]+tmp[7898]*kernel[7]+tmp[7899]*kernel[8];
				ans[7799]<=tmp[7698]*kernel[0]+tmp[7699]*kernel[1]+tmp[7798]*kernel[3]+tmp[7799]*kernel[4]+tmp[7898]*kernel[6]+tmp[7899]*kernel[7];
				ans[7800]<=tmp[7700]*kernel[1]+tmp[7701]*kernel[2]+tmp[7800]*kernel[4]+tmp[7801]*kernel[5]+tmp[7900]*kernel[7]+tmp[7901]*kernel[8];
				ans[7801]<=tmp[7700]*kernel[0]+tmp[7701]*kernel[1]+tmp[7702]*kernel[2]+tmp[7800]*kernel[3]+tmp[7801]*kernel[4]+tmp[7802]*kernel[5]+tmp[7900]*kernel[6]+tmp[7901]*kernel[7]+tmp[7902]*kernel[8];
				ans[7802]<=tmp[7701]*kernel[0]+tmp[7702]*kernel[1]+tmp[7703]*kernel[2]+tmp[7801]*kernel[3]+tmp[7802]*kernel[4]+tmp[7803]*kernel[5]+tmp[7901]*kernel[6]+tmp[7902]*kernel[7]+tmp[7903]*kernel[8];
				ans[7803]<=tmp[7702]*kernel[0]+tmp[7703]*kernel[1]+tmp[7704]*kernel[2]+tmp[7802]*kernel[3]+tmp[7803]*kernel[4]+tmp[7804]*kernel[5]+tmp[7902]*kernel[6]+tmp[7903]*kernel[7]+tmp[7904]*kernel[8];
				ans[7804]<=tmp[7703]*kernel[0]+tmp[7704]*kernel[1]+tmp[7705]*kernel[2]+tmp[7803]*kernel[3]+tmp[7804]*kernel[4]+tmp[7805]*kernel[5]+tmp[7903]*kernel[6]+tmp[7904]*kernel[7]+tmp[7905]*kernel[8];
				ans[7805]<=tmp[7704]*kernel[0]+tmp[7705]*kernel[1]+tmp[7706]*kernel[2]+tmp[7804]*kernel[3]+tmp[7805]*kernel[4]+tmp[7806]*kernel[5]+tmp[7904]*kernel[6]+tmp[7905]*kernel[7]+tmp[7906]*kernel[8];
				ans[7806]<=tmp[7705]*kernel[0]+tmp[7706]*kernel[1]+tmp[7707]*kernel[2]+tmp[7805]*kernel[3]+tmp[7806]*kernel[4]+tmp[7807]*kernel[5]+tmp[7905]*kernel[6]+tmp[7906]*kernel[7]+tmp[7907]*kernel[8];
				ans[7807]<=tmp[7706]*kernel[0]+tmp[7707]*kernel[1]+tmp[7708]*kernel[2]+tmp[7806]*kernel[3]+tmp[7807]*kernel[4]+tmp[7808]*kernel[5]+tmp[7906]*kernel[6]+tmp[7907]*kernel[7]+tmp[7908]*kernel[8];
				ans[7808]<=tmp[7707]*kernel[0]+tmp[7708]*kernel[1]+tmp[7709]*kernel[2]+tmp[7807]*kernel[3]+tmp[7808]*kernel[4]+tmp[7809]*kernel[5]+tmp[7907]*kernel[6]+tmp[7908]*kernel[7]+tmp[7909]*kernel[8];
				ans[7809]<=tmp[7708]*kernel[0]+tmp[7709]*kernel[1]+tmp[7710]*kernel[2]+tmp[7808]*kernel[3]+tmp[7809]*kernel[4]+tmp[7810]*kernel[5]+tmp[7908]*kernel[6]+tmp[7909]*kernel[7]+tmp[7910]*kernel[8];
				ans[7810]<=tmp[7709]*kernel[0]+tmp[7710]*kernel[1]+tmp[7711]*kernel[2]+tmp[7809]*kernel[3]+tmp[7810]*kernel[4]+tmp[7811]*kernel[5]+tmp[7909]*kernel[6]+tmp[7910]*kernel[7]+tmp[7911]*kernel[8];
				ans[7811]<=tmp[7710]*kernel[0]+tmp[7711]*kernel[1]+tmp[7712]*kernel[2]+tmp[7810]*kernel[3]+tmp[7811]*kernel[4]+tmp[7812]*kernel[5]+tmp[7910]*kernel[6]+tmp[7911]*kernel[7]+tmp[7912]*kernel[8];
				ans[7812]<=tmp[7711]*kernel[0]+tmp[7712]*kernel[1]+tmp[7713]*kernel[2]+tmp[7811]*kernel[3]+tmp[7812]*kernel[4]+tmp[7813]*kernel[5]+tmp[7911]*kernel[6]+tmp[7912]*kernel[7]+tmp[7913]*kernel[8];
				ans[7813]<=tmp[7712]*kernel[0]+tmp[7713]*kernel[1]+tmp[7714]*kernel[2]+tmp[7812]*kernel[3]+tmp[7813]*kernel[4]+tmp[7814]*kernel[5]+tmp[7912]*kernel[6]+tmp[7913]*kernel[7]+tmp[7914]*kernel[8];
				ans[7814]<=tmp[7713]*kernel[0]+tmp[7714]*kernel[1]+tmp[7715]*kernel[2]+tmp[7813]*kernel[3]+tmp[7814]*kernel[4]+tmp[7815]*kernel[5]+tmp[7913]*kernel[6]+tmp[7914]*kernel[7]+tmp[7915]*kernel[8];
				ans[7815]<=tmp[7714]*kernel[0]+tmp[7715]*kernel[1]+tmp[7716]*kernel[2]+tmp[7814]*kernel[3]+tmp[7815]*kernel[4]+tmp[7816]*kernel[5]+tmp[7914]*kernel[6]+tmp[7915]*kernel[7]+tmp[7916]*kernel[8];
				ans[7816]<=tmp[7715]*kernel[0]+tmp[7716]*kernel[1]+tmp[7717]*kernel[2]+tmp[7815]*kernel[3]+tmp[7816]*kernel[4]+tmp[7817]*kernel[5]+tmp[7915]*kernel[6]+tmp[7916]*kernel[7]+tmp[7917]*kernel[8];
				ans[7817]<=tmp[7716]*kernel[0]+tmp[7717]*kernel[1]+tmp[7718]*kernel[2]+tmp[7816]*kernel[3]+tmp[7817]*kernel[4]+tmp[7818]*kernel[5]+tmp[7916]*kernel[6]+tmp[7917]*kernel[7]+tmp[7918]*kernel[8];
				ans[7818]<=tmp[7717]*kernel[0]+tmp[7718]*kernel[1]+tmp[7719]*kernel[2]+tmp[7817]*kernel[3]+tmp[7818]*kernel[4]+tmp[7819]*kernel[5]+tmp[7917]*kernel[6]+tmp[7918]*kernel[7]+tmp[7919]*kernel[8];
				ans[7819]<=tmp[7718]*kernel[0]+tmp[7719]*kernel[1]+tmp[7720]*kernel[2]+tmp[7818]*kernel[3]+tmp[7819]*kernel[4]+tmp[7820]*kernel[5]+tmp[7918]*kernel[6]+tmp[7919]*kernel[7]+tmp[7920]*kernel[8];
				ans[7820]<=tmp[7719]*kernel[0]+tmp[7720]*kernel[1]+tmp[7721]*kernel[2]+tmp[7819]*kernel[3]+tmp[7820]*kernel[4]+tmp[7821]*kernel[5]+tmp[7919]*kernel[6]+tmp[7920]*kernel[7]+tmp[7921]*kernel[8];
				ans[7821]<=tmp[7720]*kernel[0]+tmp[7721]*kernel[1]+tmp[7722]*kernel[2]+tmp[7820]*kernel[3]+tmp[7821]*kernel[4]+tmp[7822]*kernel[5]+tmp[7920]*kernel[6]+tmp[7921]*kernel[7]+tmp[7922]*kernel[8];
				ans[7822]<=tmp[7721]*kernel[0]+tmp[7722]*kernel[1]+tmp[7723]*kernel[2]+tmp[7821]*kernel[3]+tmp[7822]*kernel[4]+tmp[7823]*kernel[5]+tmp[7921]*kernel[6]+tmp[7922]*kernel[7]+tmp[7923]*kernel[8];
				ans[7823]<=tmp[7722]*kernel[0]+tmp[7723]*kernel[1]+tmp[7724]*kernel[2]+tmp[7822]*kernel[3]+tmp[7823]*kernel[4]+tmp[7824]*kernel[5]+tmp[7922]*kernel[6]+tmp[7923]*kernel[7]+tmp[7924]*kernel[8];
				ans[7824]<=tmp[7723]*kernel[0]+tmp[7724]*kernel[1]+tmp[7725]*kernel[2]+tmp[7823]*kernel[3]+tmp[7824]*kernel[4]+tmp[7825]*kernel[5]+tmp[7923]*kernel[6]+tmp[7924]*kernel[7]+tmp[7925]*kernel[8];
				ans[7825]<=tmp[7724]*kernel[0]+tmp[7725]*kernel[1]+tmp[7726]*kernel[2]+tmp[7824]*kernel[3]+tmp[7825]*kernel[4]+tmp[7826]*kernel[5]+tmp[7924]*kernel[6]+tmp[7925]*kernel[7]+tmp[7926]*kernel[8];
				ans[7826]<=tmp[7725]*kernel[0]+tmp[7726]*kernel[1]+tmp[7727]*kernel[2]+tmp[7825]*kernel[3]+tmp[7826]*kernel[4]+tmp[7827]*kernel[5]+tmp[7925]*kernel[6]+tmp[7926]*kernel[7]+tmp[7927]*kernel[8];
				ans[7827]<=tmp[7726]*kernel[0]+tmp[7727]*kernel[1]+tmp[7728]*kernel[2]+tmp[7826]*kernel[3]+tmp[7827]*kernel[4]+tmp[7828]*kernel[5]+tmp[7926]*kernel[6]+tmp[7927]*kernel[7]+tmp[7928]*kernel[8];
				ans[7828]<=tmp[7727]*kernel[0]+tmp[7728]*kernel[1]+tmp[7729]*kernel[2]+tmp[7827]*kernel[3]+tmp[7828]*kernel[4]+tmp[7829]*kernel[5]+tmp[7927]*kernel[6]+tmp[7928]*kernel[7]+tmp[7929]*kernel[8];
				ans[7829]<=tmp[7728]*kernel[0]+tmp[7729]*kernel[1]+tmp[7730]*kernel[2]+tmp[7828]*kernel[3]+tmp[7829]*kernel[4]+tmp[7830]*kernel[5]+tmp[7928]*kernel[6]+tmp[7929]*kernel[7]+tmp[7930]*kernel[8];
				ans[7830]<=tmp[7729]*kernel[0]+tmp[7730]*kernel[1]+tmp[7731]*kernel[2]+tmp[7829]*kernel[3]+tmp[7830]*kernel[4]+tmp[7831]*kernel[5]+tmp[7929]*kernel[6]+tmp[7930]*kernel[7]+tmp[7931]*kernel[8];
				ans[7831]<=tmp[7730]*kernel[0]+tmp[7731]*kernel[1]+tmp[7732]*kernel[2]+tmp[7830]*kernel[3]+tmp[7831]*kernel[4]+tmp[7832]*kernel[5]+tmp[7930]*kernel[6]+tmp[7931]*kernel[7]+tmp[7932]*kernel[8];
				ans[7832]<=tmp[7731]*kernel[0]+tmp[7732]*kernel[1]+tmp[7733]*kernel[2]+tmp[7831]*kernel[3]+tmp[7832]*kernel[4]+tmp[7833]*kernel[5]+tmp[7931]*kernel[6]+tmp[7932]*kernel[7]+tmp[7933]*kernel[8];
				ans[7833]<=tmp[7732]*kernel[0]+tmp[7733]*kernel[1]+tmp[7734]*kernel[2]+tmp[7832]*kernel[3]+tmp[7833]*kernel[4]+tmp[7834]*kernel[5]+tmp[7932]*kernel[6]+tmp[7933]*kernel[7]+tmp[7934]*kernel[8];
				ans[7834]<=tmp[7733]*kernel[0]+tmp[7734]*kernel[1]+tmp[7735]*kernel[2]+tmp[7833]*kernel[3]+tmp[7834]*kernel[4]+tmp[7835]*kernel[5]+tmp[7933]*kernel[6]+tmp[7934]*kernel[7]+tmp[7935]*kernel[8];
				ans[7835]<=tmp[7734]*kernel[0]+tmp[7735]*kernel[1]+tmp[7736]*kernel[2]+tmp[7834]*kernel[3]+tmp[7835]*kernel[4]+tmp[7836]*kernel[5]+tmp[7934]*kernel[6]+tmp[7935]*kernel[7]+tmp[7936]*kernel[8];
				ans[7836]<=tmp[7735]*kernel[0]+tmp[7736]*kernel[1]+tmp[7737]*kernel[2]+tmp[7835]*kernel[3]+tmp[7836]*kernel[4]+tmp[7837]*kernel[5]+tmp[7935]*kernel[6]+tmp[7936]*kernel[7]+tmp[7937]*kernel[8];
				ans[7837]<=tmp[7736]*kernel[0]+tmp[7737]*kernel[1]+tmp[7738]*kernel[2]+tmp[7836]*kernel[3]+tmp[7837]*kernel[4]+tmp[7838]*kernel[5]+tmp[7936]*kernel[6]+tmp[7937]*kernel[7]+tmp[7938]*kernel[8];
				ans[7838]<=tmp[7737]*kernel[0]+tmp[7738]*kernel[1]+tmp[7739]*kernel[2]+tmp[7837]*kernel[3]+tmp[7838]*kernel[4]+tmp[7839]*kernel[5]+tmp[7937]*kernel[6]+tmp[7938]*kernel[7]+tmp[7939]*kernel[8];
				ans[7839]<=tmp[7738]*kernel[0]+tmp[7739]*kernel[1]+tmp[7740]*kernel[2]+tmp[7838]*kernel[3]+tmp[7839]*kernel[4]+tmp[7840]*kernel[5]+tmp[7938]*kernel[6]+tmp[7939]*kernel[7]+tmp[7940]*kernel[8];
				ans[7840]<=tmp[7739]*kernel[0]+tmp[7740]*kernel[1]+tmp[7741]*kernel[2]+tmp[7839]*kernel[3]+tmp[7840]*kernel[4]+tmp[7841]*kernel[5]+tmp[7939]*kernel[6]+tmp[7940]*kernel[7]+tmp[7941]*kernel[8];
				ans[7841]<=tmp[7740]*kernel[0]+tmp[7741]*kernel[1]+tmp[7742]*kernel[2]+tmp[7840]*kernel[3]+tmp[7841]*kernel[4]+tmp[7842]*kernel[5]+tmp[7940]*kernel[6]+tmp[7941]*kernel[7]+tmp[7942]*kernel[8];
				ans[7842]<=tmp[7741]*kernel[0]+tmp[7742]*kernel[1]+tmp[7743]*kernel[2]+tmp[7841]*kernel[3]+tmp[7842]*kernel[4]+tmp[7843]*kernel[5]+tmp[7941]*kernel[6]+tmp[7942]*kernel[7]+tmp[7943]*kernel[8];
				ans[7843]<=tmp[7742]*kernel[0]+tmp[7743]*kernel[1]+tmp[7744]*kernel[2]+tmp[7842]*kernel[3]+tmp[7843]*kernel[4]+tmp[7844]*kernel[5]+tmp[7942]*kernel[6]+tmp[7943]*kernel[7]+tmp[7944]*kernel[8];
				ans[7844]<=tmp[7743]*kernel[0]+tmp[7744]*kernel[1]+tmp[7745]*kernel[2]+tmp[7843]*kernel[3]+tmp[7844]*kernel[4]+tmp[7845]*kernel[5]+tmp[7943]*kernel[6]+tmp[7944]*kernel[7]+tmp[7945]*kernel[8];
				ans[7845]<=tmp[7744]*kernel[0]+tmp[7745]*kernel[1]+tmp[7746]*kernel[2]+tmp[7844]*kernel[3]+tmp[7845]*kernel[4]+tmp[7846]*kernel[5]+tmp[7944]*kernel[6]+tmp[7945]*kernel[7]+tmp[7946]*kernel[8];
				ans[7846]<=tmp[7745]*kernel[0]+tmp[7746]*kernel[1]+tmp[7747]*kernel[2]+tmp[7845]*kernel[3]+tmp[7846]*kernel[4]+tmp[7847]*kernel[5]+tmp[7945]*kernel[6]+tmp[7946]*kernel[7]+tmp[7947]*kernel[8];
				ans[7847]<=tmp[7746]*kernel[0]+tmp[7747]*kernel[1]+tmp[7748]*kernel[2]+tmp[7846]*kernel[3]+tmp[7847]*kernel[4]+tmp[7848]*kernel[5]+tmp[7946]*kernel[6]+tmp[7947]*kernel[7]+tmp[7948]*kernel[8];
				ans[7848]<=tmp[7747]*kernel[0]+tmp[7748]*kernel[1]+tmp[7749]*kernel[2]+tmp[7847]*kernel[3]+tmp[7848]*kernel[4]+tmp[7849]*kernel[5]+tmp[7947]*kernel[6]+tmp[7948]*kernel[7]+tmp[7949]*kernel[8];
				ans[7849]<=tmp[7748]*kernel[0]+tmp[7749]*kernel[1]+tmp[7750]*kernel[2]+tmp[7848]*kernel[3]+tmp[7849]*kernel[4]+tmp[7850]*kernel[5]+tmp[7948]*kernel[6]+tmp[7949]*kernel[7]+tmp[7950]*kernel[8];
				ans[7850]<=tmp[7749]*kernel[0]+tmp[7750]*kernel[1]+tmp[7751]*kernel[2]+tmp[7849]*kernel[3]+tmp[7850]*kernel[4]+tmp[7851]*kernel[5]+tmp[7949]*kernel[6]+tmp[7950]*kernel[7]+tmp[7951]*kernel[8];
				ans[7851]<=tmp[7750]*kernel[0]+tmp[7751]*kernel[1]+tmp[7752]*kernel[2]+tmp[7850]*kernel[3]+tmp[7851]*kernel[4]+tmp[7852]*kernel[5]+tmp[7950]*kernel[6]+tmp[7951]*kernel[7]+tmp[7952]*kernel[8];
				ans[7852]<=tmp[7751]*kernel[0]+tmp[7752]*kernel[1]+tmp[7753]*kernel[2]+tmp[7851]*kernel[3]+tmp[7852]*kernel[4]+tmp[7853]*kernel[5]+tmp[7951]*kernel[6]+tmp[7952]*kernel[7]+tmp[7953]*kernel[8];
				ans[7853]<=tmp[7752]*kernel[0]+tmp[7753]*kernel[1]+tmp[7754]*kernel[2]+tmp[7852]*kernel[3]+tmp[7853]*kernel[4]+tmp[7854]*kernel[5]+tmp[7952]*kernel[6]+tmp[7953]*kernel[7]+tmp[7954]*kernel[8];
				ans[7854]<=tmp[7753]*kernel[0]+tmp[7754]*kernel[1]+tmp[7755]*kernel[2]+tmp[7853]*kernel[3]+tmp[7854]*kernel[4]+tmp[7855]*kernel[5]+tmp[7953]*kernel[6]+tmp[7954]*kernel[7]+tmp[7955]*kernel[8];
				ans[7855]<=tmp[7754]*kernel[0]+tmp[7755]*kernel[1]+tmp[7756]*kernel[2]+tmp[7854]*kernel[3]+tmp[7855]*kernel[4]+tmp[7856]*kernel[5]+tmp[7954]*kernel[6]+tmp[7955]*kernel[7]+tmp[7956]*kernel[8];
				ans[7856]<=tmp[7755]*kernel[0]+tmp[7756]*kernel[1]+tmp[7757]*kernel[2]+tmp[7855]*kernel[3]+tmp[7856]*kernel[4]+tmp[7857]*kernel[5]+tmp[7955]*kernel[6]+tmp[7956]*kernel[7]+tmp[7957]*kernel[8];
				ans[7857]<=tmp[7756]*kernel[0]+tmp[7757]*kernel[1]+tmp[7758]*kernel[2]+tmp[7856]*kernel[3]+tmp[7857]*kernel[4]+tmp[7858]*kernel[5]+tmp[7956]*kernel[6]+tmp[7957]*kernel[7]+tmp[7958]*kernel[8];
				ans[7858]<=tmp[7757]*kernel[0]+tmp[7758]*kernel[1]+tmp[7759]*kernel[2]+tmp[7857]*kernel[3]+tmp[7858]*kernel[4]+tmp[7859]*kernel[5]+tmp[7957]*kernel[6]+tmp[7958]*kernel[7]+tmp[7959]*kernel[8];
				ans[7859]<=tmp[7758]*kernel[0]+tmp[7759]*kernel[1]+tmp[7760]*kernel[2]+tmp[7858]*kernel[3]+tmp[7859]*kernel[4]+tmp[7860]*kernel[5]+tmp[7958]*kernel[6]+tmp[7959]*kernel[7]+tmp[7960]*kernel[8];
				ans[7860]<=tmp[7759]*kernel[0]+tmp[7760]*kernel[1]+tmp[7761]*kernel[2]+tmp[7859]*kernel[3]+tmp[7860]*kernel[4]+tmp[7861]*kernel[5]+tmp[7959]*kernel[6]+tmp[7960]*kernel[7]+tmp[7961]*kernel[8];
				ans[7861]<=tmp[7760]*kernel[0]+tmp[7761]*kernel[1]+tmp[7762]*kernel[2]+tmp[7860]*kernel[3]+tmp[7861]*kernel[4]+tmp[7862]*kernel[5]+tmp[7960]*kernel[6]+tmp[7961]*kernel[7]+tmp[7962]*kernel[8];
				ans[7862]<=tmp[7761]*kernel[0]+tmp[7762]*kernel[1]+tmp[7763]*kernel[2]+tmp[7861]*kernel[3]+tmp[7862]*kernel[4]+tmp[7863]*kernel[5]+tmp[7961]*kernel[6]+tmp[7962]*kernel[7]+tmp[7963]*kernel[8];
				ans[7863]<=tmp[7762]*kernel[0]+tmp[7763]*kernel[1]+tmp[7764]*kernel[2]+tmp[7862]*kernel[3]+tmp[7863]*kernel[4]+tmp[7864]*kernel[5]+tmp[7962]*kernel[6]+tmp[7963]*kernel[7]+tmp[7964]*kernel[8];
				ans[7864]<=tmp[7763]*kernel[0]+tmp[7764]*kernel[1]+tmp[7765]*kernel[2]+tmp[7863]*kernel[3]+tmp[7864]*kernel[4]+tmp[7865]*kernel[5]+tmp[7963]*kernel[6]+tmp[7964]*kernel[7]+tmp[7965]*kernel[8];
				ans[7865]<=tmp[7764]*kernel[0]+tmp[7765]*kernel[1]+tmp[7766]*kernel[2]+tmp[7864]*kernel[3]+tmp[7865]*kernel[4]+tmp[7866]*kernel[5]+tmp[7964]*kernel[6]+tmp[7965]*kernel[7]+tmp[7966]*kernel[8];
				ans[7866]<=tmp[7765]*kernel[0]+tmp[7766]*kernel[1]+tmp[7767]*kernel[2]+tmp[7865]*kernel[3]+tmp[7866]*kernel[4]+tmp[7867]*kernel[5]+tmp[7965]*kernel[6]+tmp[7966]*kernel[7]+tmp[7967]*kernel[8];
				ans[7867]<=tmp[7766]*kernel[0]+tmp[7767]*kernel[1]+tmp[7768]*kernel[2]+tmp[7866]*kernel[3]+tmp[7867]*kernel[4]+tmp[7868]*kernel[5]+tmp[7966]*kernel[6]+tmp[7967]*kernel[7]+tmp[7968]*kernel[8];
				ans[7868]<=tmp[7767]*kernel[0]+tmp[7768]*kernel[1]+tmp[7769]*kernel[2]+tmp[7867]*kernel[3]+tmp[7868]*kernel[4]+tmp[7869]*kernel[5]+tmp[7967]*kernel[6]+tmp[7968]*kernel[7]+tmp[7969]*kernel[8];
				ans[7869]<=tmp[7768]*kernel[0]+tmp[7769]*kernel[1]+tmp[7770]*kernel[2]+tmp[7868]*kernel[3]+tmp[7869]*kernel[4]+tmp[7870]*kernel[5]+tmp[7968]*kernel[6]+tmp[7969]*kernel[7]+tmp[7970]*kernel[8];
				ans[7870]<=tmp[7769]*kernel[0]+tmp[7770]*kernel[1]+tmp[7771]*kernel[2]+tmp[7869]*kernel[3]+tmp[7870]*kernel[4]+tmp[7871]*kernel[5]+tmp[7969]*kernel[6]+tmp[7970]*kernel[7]+tmp[7971]*kernel[8];
				ans[7871]<=tmp[7770]*kernel[0]+tmp[7771]*kernel[1]+tmp[7772]*kernel[2]+tmp[7870]*kernel[3]+tmp[7871]*kernel[4]+tmp[7872]*kernel[5]+tmp[7970]*kernel[6]+tmp[7971]*kernel[7]+tmp[7972]*kernel[8];
				ans[7872]<=tmp[7771]*kernel[0]+tmp[7772]*kernel[1]+tmp[7773]*kernel[2]+tmp[7871]*kernel[3]+tmp[7872]*kernel[4]+tmp[7873]*kernel[5]+tmp[7971]*kernel[6]+tmp[7972]*kernel[7]+tmp[7973]*kernel[8];
				ans[7873]<=tmp[7772]*kernel[0]+tmp[7773]*kernel[1]+tmp[7774]*kernel[2]+tmp[7872]*kernel[3]+tmp[7873]*kernel[4]+tmp[7874]*kernel[5]+tmp[7972]*kernel[6]+tmp[7973]*kernel[7]+tmp[7974]*kernel[8];
				ans[7874]<=tmp[7773]*kernel[0]+tmp[7774]*kernel[1]+tmp[7775]*kernel[2]+tmp[7873]*kernel[3]+tmp[7874]*kernel[4]+tmp[7875]*kernel[5]+tmp[7973]*kernel[6]+tmp[7974]*kernel[7]+tmp[7975]*kernel[8];
				ans[7875]<=tmp[7774]*kernel[0]+tmp[7775]*kernel[1]+tmp[7776]*kernel[2]+tmp[7874]*kernel[3]+tmp[7875]*kernel[4]+tmp[7876]*kernel[5]+tmp[7974]*kernel[6]+tmp[7975]*kernel[7]+tmp[7976]*kernel[8];
				ans[7876]<=tmp[7775]*kernel[0]+tmp[7776]*kernel[1]+tmp[7777]*kernel[2]+tmp[7875]*kernel[3]+tmp[7876]*kernel[4]+tmp[7877]*kernel[5]+tmp[7975]*kernel[6]+tmp[7976]*kernel[7]+tmp[7977]*kernel[8];
				ans[7877]<=tmp[7776]*kernel[0]+tmp[7777]*kernel[1]+tmp[7778]*kernel[2]+tmp[7876]*kernel[3]+tmp[7877]*kernel[4]+tmp[7878]*kernel[5]+tmp[7976]*kernel[6]+tmp[7977]*kernel[7]+tmp[7978]*kernel[8];
				ans[7878]<=tmp[7777]*kernel[0]+tmp[7778]*kernel[1]+tmp[7779]*kernel[2]+tmp[7877]*kernel[3]+tmp[7878]*kernel[4]+tmp[7879]*kernel[5]+tmp[7977]*kernel[6]+tmp[7978]*kernel[7]+tmp[7979]*kernel[8];
				ans[7879]<=tmp[7778]*kernel[0]+tmp[7779]*kernel[1]+tmp[7780]*kernel[2]+tmp[7878]*kernel[3]+tmp[7879]*kernel[4]+tmp[7880]*kernel[5]+tmp[7978]*kernel[6]+tmp[7979]*kernel[7]+tmp[7980]*kernel[8];
				ans[7880]<=tmp[7779]*kernel[0]+tmp[7780]*kernel[1]+tmp[7781]*kernel[2]+tmp[7879]*kernel[3]+tmp[7880]*kernel[4]+tmp[7881]*kernel[5]+tmp[7979]*kernel[6]+tmp[7980]*kernel[7]+tmp[7981]*kernel[8];
				ans[7881]<=tmp[7780]*kernel[0]+tmp[7781]*kernel[1]+tmp[7782]*kernel[2]+tmp[7880]*kernel[3]+tmp[7881]*kernel[4]+tmp[7882]*kernel[5]+tmp[7980]*kernel[6]+tmp[7981]*kernel[7]+tmp[7982]*kernel[8];
				ans[7882]<=tmp[7781]*kernel[0]+tmp[7782]*kernel[1]+tmp[7783]*kernel[2]+tmp[7881]*kernel[3]+tmp[7882]*kernel[4]+tmp[7883]*kernel[5]+tmp[7981]*kernel[6]+tmp[7982]*kernel[7]+tmp[7983]*kernel[8];
				ans[7883]<=tmp[7782]*kernel[0]+tmp[7783]*kernel[1]+tmp[7784]*kernel[2]+tmp[7882]*kernel[3]+tmp[7883]*kernel[4]+tmp[7884]*kernel[5]+tmp[7982]*kernel[6]+tmp[7983]*kernel[7]+tmp[7984]*kernel[8];
				ans[7884]<=tmp[7783]*kernel[0]+tmp[7784]*kernel[1]+tmp[7785]*kernel[2]+tmp[7883]*kernel[3]+tmp[7884]*kernel[4]+tmp[7885]*kernel[5]+tmp[7983]*kernel[6]+tmp[7984]*kernel[7]+tmp[7985]*kernel[8];
				ans[7885]<=tmp[7784]*kernel[0]+tmp[7785]*kernel[1]+tmp[7786]*kernel[2]+tmp[7884]*kernel[3]+tmp[7885]*kernel[4]+tmp[7886]*kernel[5]+tmp[7984]*kernel[6]+tmp[7985]*kernel[7]+tmp[7986]*kernel[8];
				ans[7886]<=tmp[7785]*kernel[0]+tmp[7786]*kernel[1]+tmp[7787]*kernel[2]+tmp[7885]*kernel[3]+tmp[7886]*kernel[4]+tmp[7887]*kernel[5]+tmp[7985]*kernel[6]+tmp[7986]*kernel[7]+tmp[7987]*kernel[8];
				ans[7887]<=tmp[7786]*kernel[0]+tmp[7787]*kernel[1]+tmp[7788]*kernel[2]+tmp[7886]*kernel[3]+tmp[7887]*kernel[4]+tmp[7888]*kernel[5]+tmp[7986]*kernel[6]+tmp[7987]*kernel[7]+tmp[7988]*kernel[8];
				ans[7888]<=tmp[7787]*kernel[0]+tmp[7788]*kernel[1]+tmp[7789]*kernel[2]+tmp[7887]*kernel[3]+tmp[7888]*kernel[4]+tmp[7889]*kernel[5]+tmp[7987]*kernel[6]+tmp[7988]*kernel[7]+tmp[7989]*kernel[8];
				ans[7889]<=tmp[7788]*kernel[0]+tmp[7789]*kernel[1]+tmp[7790]*kernel[2]+tmp[7888]*kernel[3]+tmp[7889]*kernel[4]+tmp[7890]*kernel[5]+tmp[7988]*kernel[6]+tmp[7989]*kernel[7]+tmp[7990]*kernel[8];
				ans[7890]<=tmp[7789]*kernel[0]+tmp[7790]*kernel[1]+tmp[7791]*kernel[2]+tmp[7889]*kernel[3]+tmp[7890]*kernel[4]+tmp[7891]*kernel[5]+tmp[7989]*kernel[6]+tmp[7990]*kernel[7]+tmp[7991]*kernel[8];
				ans[7891]<=tmp[7790]*kernel[0]+tmp[7791]*kernel[1]+tmp[7792]*kernel[2]+tmp[7890]*kernel[3]+tmp[7891]*kernel[4]+tmp[7892]*kernel[5]+tmp[7990]*kernel[6]+tmp[7991]*kernel[7]+tmp[7992]*kernel[8];
				ans[7892]<=tmp[7791]*kernel[0]+tmp[7792]*kernel[1]+tmp[7793]*kernel[2]+tmp[7891]*kernel[3]+tmp[7892]*kernel[4]+tmp[7893]*kernel[5]+tmp[7991]*kernel[6]+tmp[7992]*kernel[7]+tmp[7993]*kernel[8];
				ans[7893]<=tmp[7792]*kernel[0]+tmp[7793]*kernel[1]+tmp[7794]*kernel[2]+tmp[7892]*kernel[3]+tmp[7893]*kernel[4]+tmp[7894]*kernel[5]+tmp[7992]*kernel[6]+tmp[7993]*kernel[7]+tmp[7994]*kernel[8];
				ans[7894]<=tmp[7793]*kernel[0]+tmp[7794]*kernel[1]+tmp[7795]*kernel[2]+tmp[7893]*kernel[3]+tmp[7894]*kernel[4]+tmp[7895]*kernel[5]+tmp[7993]*kernel[6]+tmp[7994]*kernel[7]+tmp[7995]*kernel[8];
				ans[7895]<=tmp[7794]*kernel[0]+tmp[7795]*kernel[1]+tmp[7796]*kernel[2]+tmp[7894]*kernel[3]+tmp[7895]*kernel[4]+tmp[7896]*kernel[5]+tmp[7994]*kernel[6]+tmp[7995]*kernel[7]+tmp[7996]*kernel[8];
				ans[7896]<=tmp[7795]*kernel[0]+tmp[7796]*kernel[1]+tmp[7797]*kernel[2]+tmp[7895]*kernel[3]+tmp[7896]*kernel[4]+tmp[7897]*kernel[5]+tmp[7995]*kernel[6]+tmp[7996]*kernel[7]+tmp[7997]*kernel[8];
				ans[7897]<=tmp[7796]*kernel[0]+tmp[7797]*kernel[1]+tmp[7798]*kernel[2]+tmp[7896]*kernel[3]+tmp[7897]*kernel[4]+tmp[7898]*kernel[5]+tmp[7996]*kernel[6]+tmp[7997]*kernel[7]+tmp[7998]*kernel[8];
				ans[7898]<=tmp[7797]*kernel[0]+tmp[7798]*kernel[1]+tmp[7799]*kernel[2]+tmp[7897]*kernel[3]+tmp[7898]*kernel[4]+tmp[7899]*kernel[5]+tmp[7997]*kernel[6]+tmp[7998]*kernel[7]+tmp[7999]*kernel[8];
				ans[7899]<=tmp[7798]*kernel[0]+tmp[7799]*kernel[1]+tmp[7898]*kernel[3]+tmp[7899]*kernel[4]+tmp[7998]*kernel[6]+tmp[7999]*kernel[7];
				ans[7900]<=tmp[7800]*kernel[1]+tmp[7801]*kernel[2]+tmp[7900]*kernel[4]+tmp[7901]*kernel[5]+tmp[8000]*kernel[7]+tmp[8001]*kernel[8];
				ans[7901]<=tmp[7800]*kernel[0]+tmp[7801]*kernel[1]+tmp[7802]*kernel[2]+tmp[7900]*kernel[3]+tmp[7901]*kernel[4]+tmp[7902]*kernel[5]+tmp[8000]*kernel[6]+tmp[8001]*kernel[7]+tmp[8002]*kernel[8];
				ans[7902]<=tmp[7801]*kernel[0]+tmp[7802]*kernel[1]+tmp[7803]*kernel[2]+tmp[7901]*kernel[3]+tmp[7902]*kernel[4]+tmp[7903]*kernel[5]+tmp[8001]*kernel[6]+tmp[8002]*kernel[7]+tmp[8003]*kernel[8];
				ans[7903]<=tmp[7802]*kernel[0]+tmp[7803]*kernel[1]+tmp[7804]*kernel[2]+tmp[7902]*kernel[3]+tmp[7903]*kernel[4]+tmp[7904]*kernel[5]+tmp[8002]*kernel[6]+tmp[8003]*kernel[7]+tmp[8004]*kernel[8];
				ans[7904]<=tmp[7803]*kernel[0]+tmp[7804]*kernel[1]+tmp[7805]*kernel[2]+tmp[7903]*kernel[3]+tmp[7904]*kernel[4]+tmp[7905]*kernel[5]+tmp[8003]*kernel[6]+tmp[8004]*kernel[7]+tmp[8005]*kernel[8];
				ans[7905]<=tmp[7804]*kernel[0]+tmp[7805]*kernel[1]+tmp[7806]*kernel[2]+tmp[7904]*kernel[3]+tmp[7905]*kernel[4]+tmp[7906]*kernel[5]+tmp[8004]*kernel[6]+tmp[8005]*kernel[7]+tmp[8006]*kernel[8];
				ans[7906]<=tmp[7805]*kernel[0]+tmp[7806]*kernel[1]+tmp[7807]*kernel[2]+tmp[7905]*kernel[3]+tmp[7906]*kernel[4]+tmp[7907]*kernel[5]+tmp[8005]*kernel[6]+tmp[8006]*kernel[7]+tmp[8007]*kernel[8];
				ans[7907]<=tmp[7806]*kernel[0]+tmp[7807]*kernel[1]+tmp[7808]*kernel[2]+tmp[7906]*kernel[3]+tmp[7907]*kernel[4]+tmp[7908]*kernel[5]+tmp[8006]*kernel[6]+tmp[8007]*kernel[7]+tmp[8008]*kernel[8];
				ans[7908]<=tmp[7807]*kernel[0]+tmp[7808]*kernel[1]+tmp[7809]*kernel[2]+tmp[7907]*kernel[3]+tmp[7908]*kernel[4]+tmp[7909]*kernel[5]+tmp[8007]*kernel[6]+tmp[8008]*kernel[7]+tmp[8009]*kernel[8];
				ans[7909]<=tmp[7808]*kernel[0]+tmp[7809]*kernel[1]+tmp[7810]*kernel[2]+tmp[7908]*kernel[3]+tmp[7909]*kernel[4]+tmp[7910]*kernel[5]+tmp[8008]*kernel[6]+tmp[8009]*kernel[7]+tmp[8010]*kernel[8];
				ans[7910]<=tmp[7809]*kernel[0]+tmp[7810]*kernel[1]+tmp[7811]*kernel[2]+tmp[7909]*kernel[3]+tmp[7910]*kernel[4]+tmp[7911]*kernel[5]+tmp[8009]*kernel[6]+tmp[8010]*kernel[7]+tmp[8011]*kernel[8];
				ans[7911]<=tmp[7810]*kernel[0]+tmp[7811]*kernel[1]+tmp[7812]*kernel[2]+tmp[7910]*kernel[3]+tmp[7911]*kernel[4]+tmp[7912]*kernel[5]+tmp[8010]*kernel[6]+tmp[8011]*kernel[7]+tmp[8012]*kernel[8];
				ans[7912]<=tmp[7811]*kernel[0]+tmp[7812]*kernel[1]+tmp[7813]*kernel[2]+tmp[7911]*kernel[3]+tmp[7912]*kernel[4]+tmp[7913]*kernel[5]+tmp[8011]*kernel[6]+tmp[8012]*kernel[7]+tmp[8013]*kernel[8];
				ans[7913]<=tmp[7812]*kernel[0]+tmp[7813]*kernel[1]+tmp[7814]*kernel[2]+tmp[7912]*kernel[3]+tmp[7913]*kernel[4]+tmp[7914]*kernel[5]+tmp[8012]*kernel[6]+tmp[8013]*kernel[7]+tmp[8014]*kernel[8];
				ans[7914]<=tmp[7813]*kernel[0]+tmp[7814]*kernel[1]+tmp[7815]*kernel[2]+tmp[7913]*kernel[3]+tmp[7914]*kernel[4]+tmp[7915]*kernel[5]+tmp[8013]*kernel[6]+tmp[8014]*kernel[7]+tmp[8015]*kernel[8];
				ans[7915]<=tmp[7814]*kernel[0]+tmp[7815]*kernel[1]+tmp[7816]*kernel[2]+tmp[7914]*kernel[3]+tmp[7915]*kernel[4]+tmp[7916]*kernel[5]+tmp[8014]*kernel[6]+tmp[8015]*kernel[7]+tmp[8016]*kernel[8];
				ans[7916]<=tmp[7815]*kernel[0]+tmp[7816]*kernel[1]+tmp[7817]*kernel[2]+tmp[7915]*kernel[3]+tmp[7916]*kernel[4]+tmp[7917]*kernel[5]+tmp[8015]*kernel[6]+tmp[8016]*kernel[7]+tmp[8017]*kernel[8];
				ans[7917]<=tmp[7816]*kernel[0]+tmp[7817]*kernel[1]+tmp[7818]*kernel[2]+tmp[7916]*kernel[3]+tmp[7917]*kernel[4]+tmp[7918]*kernel[5]+tmp[8016]*kernel[6]+tmp[8017]*kernel[7]+tmp[8018]*kernel[8];
				ans[7918]<=tmp[7817]*kernel[0]+tmp[7818]*kernel[1]+tmp[7819]*kernel[2]+tmp[7917]*kernel[3]+tmp[7918]*kernel[4]+tmp[7919]*kernel[5]+tmp[8017]*kernel[6]+tmp[8018]*kernel[7]+tmp[8019]*kernel[8];
				ans[7919]<=tmp[7818]*kernel[0]+tmp[7819]*kernel[1]+tmp[7820]*kernel[2]+tmp[7918]*kernel[3]+tmp[7919]*kernel[4]+tmp[7920]*kernel[5]+tmp[8018]*kernel[6]+tmp[8019]*kernel[7]+tmp[8020]*kernel[8];
				ans[7920]<=tmp[7819]*kernel[0]+tmp[7820]*kernel[1]+tmp[7821]*kernel[2]+tmp[7919]*kernel[3]+tmp[7920]*kernel[4]+tmp[7921]*kernel[5]+tmp[8019]*kernel[6]+tmp[8020]*kernel[7]+tmp[8021]*kernel[8];
				ans[7921]<=tmp[7820]*kernel[0]+tmp[7821]*kernel[1]+tmp[7822]*kernel[2]+tmp[7920]*kernel[3]+tmp[7921]*kernel[4]+tmp[7922]*kernel[5]+tmp[8020]*kernel[6]+tmp[8021]*kernel[7]+tmp[8022]*kernel[8];
				ans[7922]<=tmp[7821]*kernel[0]+tmp[7822]*kernel[1]+tmp[7823]*kernel[2]+tmp[7921]*kernel[3]+tmp[7922]*kernel[4]+tmp[7923]*kernel[5]+tmp[8021]*kernel[6]+tmp[8022]*kernel[7]+tmp[8023]*kernel[8];
				ans[7923]<=tmp[7822]*kernel[0]+tmp[7823]*kernel[1]+tmp[7824]*kernel[2]+tmp[7922]*kernel[3]+tmp[7923]*kernel[4]+tmp[7924]*kernel[5]+tmp[8022]*kernel[6]+tmp[8023]*kernel[7]+tmp[8024]*kernel[8];
				ans[7924]<=tmp[7823]*kernel[0]+tmp[7824]*kernel[1]+tmp[7825]*kernel[2]+tmp[7923]*kernel[3]+tmp[7924]*kernel[4]+tmp[7925]*kernel[5]+tmp[8023]*kernel[6]+tmp[8024]*kernel[7]+tmp[8025]*kernel[8];
				ans[7925]<=tmp[7824]*kernel[0]+tmp[7825]*kernel[1]+tmp[7826]*kernel[2]+tmp[7924]*kernel[3]+tmp[7925]*kernel[4]+tmp[7926]*kernel[5]+tmp[8024]*kernel[6]+tmp[8025]*kernel[7]+tmp[8026]*kernel[8];
				ans[7926]<=tmp[7825]*kernel[0]+tmp[7826]*kernel[1]+tmp[7827]*kernel[2]+tmp[7925]*kernel[3]+tmp[7926]*kernel[4]+tmp[7927]*kernel[5]+tmp[8025]*kernel[6]+tmp[8026]*kernel[7]+tmp[8027]*kernel[8];
				ans[7927]<=tmp[7826]*kernel[0]+tmp[7827]*kernel[1]+tmp[7828]*kernel[2]+tmp[7926]*kernel[3]+tmp[7927]*kernel[4]+tmp[7928]*kernel[5]+tmp[8026]*kernel[6]+tmp[8027]*kernel[7]+tmp[8028]*kernel[8];
				ans[7928]<=tmp[7827]*kernel[0]+tmp[7828]*kernel[1]+tmp[7829]*kernel[2]+tmp[7927]*kernel[3]+tmp[7928]*kernel[4]+tmp[7929]*kernel[5]+tmp[8027]*kernel[6]+tmp[8028]*kernel[7]+tmp[8029]*kernel[8];
				ans[7929]<=tmp[7828]*kernel[0]+tmp[7829]*kernel[1]+tmp[7830]*kernel[2]+tmp[7928]*kernel[3]+tmp[7929]*kernel[4]+tmp[7930]*kernel[5]+tmp[8028]*kernel[6]+tmp[8029]*kernel[7]+tmp[8030]*kernel[8];
				ans[7930]<=tmp[7829]*kernel[0]+tmp[7830]*kernel[1]+tmp[7831]*kernel[2]+tmp[7929]*kernel[3]+tmp[7930]*kernel[4]+tmp[7931]*kernel[5]+tmp[8029]*kernel[6]+tmp[8030]*kernel[7]+tmp[8031]*kernel[8];
				ans[7931]<=tmp[7830]*kernel[0]+tmp[7831]*kernel[1]+tmp[7832]*kernel[2]+tmp[7930]*kernel[3]+tmp[7931]*kernel[4]+tmp[7932]*kernel[5]+tmp[8030]*kernel[6]+tmp[8031]*kernel[7]+tmp[8032]*kernel[8];
				ans[7932]<=tmp[7831]*kernel[0]+tmp[7832]*kernel[1]+tmp[7833]*kernel[2]+tmp[7931]*kernel[3]+tmp[7932]*kernel[4]+tmp[7933]*kernel[5]+tmp[8031]*kernel[6]+tmp[8032]*kernel[7]+tmp[8033]*kernel[8];
				ans[7933]<=tmp[7832]*kernel[0]+tmp[7833]*kernel[1]+tmp[7834]*kernel[2]+tmp[7932]*kernel[3]+tmp[7933]*kernel[4]+tmp[7934]*kernel[5]+tmp[8032]*kernel[6]+tmp[8033]*kernel[7]+tmp[8034]*kernel[8];
				ans[7934]<=tmp[7833]*kernel[0]+tmp[7834]*kernel[1]+tmp[7835]*kernel[2]+tmp[7933]*kernel[3]+tmp[7934]*kernel[4]+tmp[7935]*kernel[5]+tmp[8033]*kernel[6]+tmp[8034]*kernel[7]+tmp[8035]*kernel[8];
				ans[7935]<=tmp[7834]*kernel[0]+tmp[7835]*kernel[1]+tmp[7836]*kernel[2]+tmp[7934]*kernel[3]+tmp[7935]*kernel[4]+tmp[7936]*kernel[5]+tmp[8034]*kernel[6]+tmp[8035]*kernel[7]+tmp[8036]*kernel[8];
				ans[7936]<=tmp[7835]*kernel[0]+tmp[7836]*kernel[1]+tmp[7837]*kernel[2]+tmp[7935]*kernel[3]+tmp[7936]*kernel[4]+tmp[7937]*kernel[5]+tmp[8035]*kernel[6]+tmp[8036]*kernel[7]+tmp[8037]*kernel[8];
				ans[7937]<=tmp[7836]*kernel[0]+tmp[7837]*kernel[1]+tmp[7838]*kernel[2]+tmp[7936]*kernel[3]+tmp[7937]*kernel[4]+tmp[7938]*kernel[5]+tmp[8036]*kernel[6]+tmp[8037]*kernel[7]+tmp[8038]*kernel[8];
				ans[7938]<=tmp[7837]*kernel[0]+tmp[7838]*kernel[1]+tmp[7839]*kernel[2]+tmp[7937]*kernel[3]+tmp[7938]*kernel[4]+tmp[7939]*kernel[5]+tmp[8037]*kernel[6]+tmp[8038]*kernel[7]+tmp[8039]*kernel[8];
				ans[7939]<=tmp[7838]*kernel[0]+tmp[7839]*kernel[1]+tmp[7840]*kernel[2]+tmp[7938]*kernel[3]+tmp[7939]*kernel[4]+tmp[7940]*kernel[5]+tmp[8038]*kernel[6]+tmp[8039]*kernel[7]+tmp[8040]*kernel[8];
				ans[7940]<=tmp[7839]*kernel[0]+tmp[7840]*kernel[1]+tmp[7841]*kernel[2]+tmp[7939]*kernel[3]+tmp[7940]*kernel[4]+tmp[7941]*kernel[5]+tmp[8039]*kernel[6]+tmp[8040]*kernel[7]+tmp[8041]*kernel[8];
				ans[7941]<=tmp[7840]*kernel[0]+tmp[7841]*kernel[1]+tmp[7842]*kernel[2]+tmp[7940]*kernel[3]+tmp[7941]*kernel[4]+tmp[7942]*kernel[5]+tmp[8040]*kernel[6]+tmp[8041]*kernel[7]+tmp[8042]*kernel[8];
				ans[7942]<=tmp[7841]*kernel[0]+tmp[7842]*kernel[1]+tmp[7843]*kernel[2]+tmp[7941]*kernel[3]+tmp[7942]*kernel[4]+tmp[7943]*kernel[5]+tmp[8041]*kernel[6]+tmp[8042]*kernel[7]+tmp[8043]*kernel[8];
				ans[7943]<=tmp[7842]*kernel[0]+tmp[7843]*kernel[1]+tmp[7844]*kernel[2]+tmp[7942]*kernel[3]+tmp[7943]*kernel[4]+tmp[7944]*kernel[5]+tmp[8042]*kernel[6]+tmp[8043]*kernel[7]+tmp[8044]*kernel[8];
				ans[7944]<=tmp[7843]*kernel[0]+tmp[7844]*kernel[1]+tmp[7845]*kernel[2]+tmp[7943]*kernel[3]+tmp[7944]*kernel[4]+tmp[7945]*kernel[5]+tmp[8043]*kernel[6]+tmp[8044]*kernel[7]+tmp[8045]*kernel[8];
				ans[7945]<=tmp[7844]*kernel[0]+tmp[7845]*kernel[1]+tmp[7846]*kernel[2]+tmp[7944]*kernel[3]+tmp[7945]*kernel[4]+tmp[7946]*kernel[5]+tmp[8044]*kernel[6]+tmp[8045]*kernel[7]+tmp[8046]*kernel[8];
				ans[7946]<=tmp[7845]*kernel[0]+tmp[7846]*kernel[1]+tmp[7847]*kernel[2]+tmp[7945]*kernel[3]+tmp[7946]*kernel[4]+tmp[7947]*kernel[5]+tmp[8045]*kernel[6]+tmp[8046]*kernel[7]+tmp[8047]*kernel[8];
				ans[7947]<=tmp[7846]*kernel[0]+tmp[7847]*kernel[1]+tmp[7848]*kernel[2]+tmp[7946]*kernel[3]+tmp[7947]*kernel[4]+tmp[7948]*kernel[5]+tmp[8046]*kernel[6]+tmp[8047]*kernel[7]+tmp[8048]*kernel[8];
				ans[7948]<=tmp[7847]*kernel[0]+tmp[7848]*kernel[1]+tmp[7849]*kernel[2]+tmp[7947]*kernel[3]+tmp[7948]*kernel[4]+tmp[7949]*kernel[5]+tmp[8047]*kernel[6]+tmp[8048]*kernel[7]+tmp[8049]*kernel[8];
				ans[7949]<=tmp[7848]*kernel[0]+tmp[7849]*kernel[1]+tmp[7850]*kernel[2]+tmp[7948]*kernel[3]+tmp[7949]*kernel[4]+tmp[7950]*kernel[5]+tmp[8048]*kernel[6]+tmp[8049]*kernel[7]+tmp[8050]*kernel[8];
				ans[7950]<=tmp[7849]*kernel[0]+tmp[7850]*kernel[1]+tmp[7851]*kernel[2]+tmp[7949]*kernel[3]+tmp[7950]*kernel[4]+tmp[7951]*kernel[5]+tmp[8049]*kernel[6]+tmp[8050]*kernel[7]+tmp[8051]*kernel[8];
				ans[7951]<=tmp[7850]*kernel[0]+tmp[7851]*kernel[1]+tmp[7852]*kernel[2]+tmp[7950]*kernel[3]+tmp[7951]*kernel[4]+tmp[7952]*kernel[5]+tmp[8050]*kernel[6]+tmp[8051]*kernel[7]+tmp[8052]*kernel[8];
				ans[7952]<=tmp[7851]*kernel[0]+tmp[7852]*kernel[1]+tmp[7853]*kernel[2]+tmp[7951]*kernel[3]+tmp[7952]*kernel[4]+tmp[7953]*kernel[5]+tmp[8051]*kernel[6]+tmp[8052]*kernel[7]+tmp[8053]*kernel[8];
				ans[7953]<=tmp[7852]*kernel[0]+tmp[7853]*kernel[1]+tmp[7854]*kernel[2]+tmp[7952]*kernel[3]+tmp[7953]*kernel[4]+tmp[7954]*kernel[5]+tmp[8052]*kernel[6]+tmp[8053]*kernel[7]+tmp[8054]*kernel[8];
				ans[7954]<=tmp[7853]*kernel[0]+tmp[7854]*kernel[1]+tmp[7855]*kernel[2]+tmp[7953]*kernel[3]+tmp[7954]*kernel[4]+tmp[7955]*kernel[5]+tmp[8053]*kernel[6]+tmp[8054]*kernel[7]+tmp[8055]*kernel[8];
				ans[7955]<=tmp[7854]*kernel[0]+tmp[7855]*kernel[1]+tmp[7856]*kernel[2]+tmp[7954]*kernel[3]+tmp[7955]*kernel[4]+tmp[7956]*kernel[5]+tmp[8054]*kernel[6]+tmp[8055]*kernel[7]+tmp[8056]*kernel[8];
				ans[7956]<=tmp[7855]*kernel[0]+tmp[7856]*kernel[1]+tmp[7857]*kernel[2]+tmp[7955]*kernel[3]+tmp[7956]*kernel[4]+tmp[7957]*kernel[5]+tmp[8055]*kernel[6]+tmp[8056]*kernel[7]+tmp[8057]*kernel[8];
				ans[7957]<=tmp[7856]*kernel[0]+tmp[7857]*kernel[1]+tmp[7858]*kernel[2]+tmp[7956]*kernel[3]+tmp[7957]*kernel[4]+tmp[7958]*kernel[5]+tmp[8056]*kernel[6]+tmp[8057]*kernel[7]+tmp[8058]*kernel[8];
				ans[7958]<=tmp[7857]*kernel[0]+tmp[7858]*kernel[1]+tmp[7859]*kernel[2]+tmp[7957]*kernel[3]+tmp[7958]*kernel[4]+tmp[7959]*kernel[5]+tmp[8057]*kernel[6]+tmp[8058]*kernel[7]+tmp[8059]*kernel[8];
				ans[7959]<=tmp[7858]*kernel[0]+tmp[7859]*kernel[1]+tmp[7860]*kernel[2]+tmp[7958]*kernel[3]+tmp[7959]*kernel[4]+tmp[7960]*kernel[5]+tmp[8058]*kernel[6]+tmp[8059]*kernel[7]+tmp[8060]*kernel[8];
				ans[7960]<=tmp[7859]*kernel[0]+tmp[7860]*kernel[1]+tmp[7861]*kernel[2]+tmp[7959]*kernel[3]+tmp[7960]*kernel[4]+tmp[7961]*kernel[5]+tmp[8059]*kernel[6]+tmp[8060]*kernel[7]+tmp[8061]*kernel[8];
				ans[7961]<=tmp[7860]*kernel[0]+tmp[7861]*kernel[1]+tmp[7862]*kernel[2]+tmp[7960]*kernel[3]+tmp[7961]*kernel[4]+tmp[7962]*kernel[5]+tmp[8060]*kernel[6]+tmp[8061]*kernel[7]+tmp[8062]*kernel[8];
				ans[7962]<=tmp[7861]*kernel[0]+tmp[7862]*kernel[1]+tmp[7863]*kernel[2]+tmp[7961]*kernel[3]+tmp[7962]*kernel[4]+tmp[7963]*kernel[5]+tmp[8061]*kernel[6]+tmp[8062]*kernel[7]+tmp[8063]*kernel[8];
				ans[7963]<=tmp[7862]*kernel[0]+tmp[7863]*kernel[1]+tmp[7864]*kernel[2]+tmp[7962]*kernel[3]+tmp[7963]*kernel[4]+tmp[7964]*kernel[5]+tmp[8062]*kernel[6]+tmp[8063]*kernel[7]+tmp[8064]*kernel[8];
				ans[7964]<=tmp[7863]*kernel[0]+tmp[7864]*kernel[1]+tmp[7865]*kernel[2]+tmp[7963]*kernel[3]+tmp[7964]*kernel[4]+tmp[7965]*kernel[5]+tmp[8063]*kernel[6]+tmp[8064]*kernel[7]+tmp[8065]*kernel[8];
				ans[7965]<=tmp[7864]*kernel[0]+tmp[7865]*kernel[1]+tmp[7866]*kernel[2]+tmp[7964]*kernel[3]+tmp[7965]*kernel[4]+tmp[7966]*kernel[5]+tmp[8064]*kernel[6]+tmp[8065]*kernel[7]+tmp[8066]*kernel[8];
				ans[7966]<=tmp[7865]*kernel[0]+tmp[7866]*kernel[1]+tmp[7867]*kernel[2]+tmp[7965]*kernel[3]+tmp[7966]*kernel[4]+tmp[7967]*kernel[5]+tmp[8065]*kernel[6]+tmp[8066]*kernel[7]+tmp[8067]*kernel[8];
				ans[7967]<=tmp[7866]*kernel[0]+tmp[7867]*kernel[1]+tmp[7868]*kernel[2]+tmp[7966]*kernel[3]+tmp[7967]*kernel[4]+tmp[7968]*kernel[5]+tmp[8066]*kernel[6]+tmp[8067]*kernel[7]+tmp[8068]*kernel[8];
				ans[7968]<=tmp[7867]*kernel[0]+tmp[7868]*kernel[1]+tmp[7869]*kernel[2]+tmp[7967]*kernel[3]+tmp[7968]*kernel[4]+tmp[7969]*kernel[5]+tmp[8067]*kernel[6]+tmp[8068]*kernel[7]+tmp[8069]*kernel[8];
				ans[7969]<=tmp[7868]*kernel[0]+tmp[7869]*kernel[1]+tmp[7870]*kernel[2]+tmp[7968]*kernel[3]+tmp[7969]*kernel[4]+tmp[7970]*kernel[5]+tmp[8068]*kernel[6]+tmp[8069]*kernel[7]+tmp[8070]*kernel[8];
				ans[7970]<=tmp[7869]*kernel[0]+tmp[7870]*kernel[1]+tmp[7871]*kernel[2]+tmp[7969]*kernel[3]+tmp[7970]*kernel[4]+tmp[7971]*kernel[5]+tmp[8069]*kernel[6]+tmp[8070]*kernel[7]+tmp[8071]*kernel[8];
				ans[7971]<=tmp[7870]*kernel[0]+tmp[7871]*kernel[1]+tmp[7872]*kernel[2]+tmp[7970]*kernel[3]+tmp[7971]*kernel[4]+tmp[7972]*kernel[5]+tmp[8070]*kernel[6]+tmp[8071]*kernel[7]+tmp[8072]*kernel[8];
				ans[7972]<=tmp[7871]*kernel[0]+tmp[7872]*kernel[1]+tmp[7873]*kernel[2]+tmp[7971]*kernel[3]+tmp[7972]*kernel[4]+tmp[7973]*kernel[5]+tmp[8071]*kernel[6]+tmp[8072]*kernel[7]+tmp[8073]*kernel[8];
				ans[7973]<=tmp[7872]*kernel[0]+tmp[7873]*kernel[1]+tmp[7874]*kernel[2]+tmp[7972]*kernel[3]+tmp[7973]*kernel[4]+tmp[7974]*kernel[5]+tmp[8072]*kernel[6]+tmp[8073]*kernel[7]+tmp[8074]*kernel[8];
				ans[7974]<=tmp[7873]*kernel[0]+tmp[7874]*kernel[1]+tmp[7875]*kernel[2]+tmp[7973]*kernel[3]+tmp[7974]*kernel[4]+tmp[7975]*kernel[5]+tmp[8073]*kernel[6]+tmp[8074]*kernel[7]+tmp[8075]*kernel[8];
				ans[7975]<=tmp[7874]*kernel[0]+tmp[7875]*kernel[1]+tmp[7876]*kernel[2]+tmp[7974]*kernel[3]+tmp[7975]*kernel[4]+tmp[7976]*kernel[5]+tmp[8074]*kernel[6]+tmp[8075]*kernel[7]+tmp[8076]*kernel[8];
				ans[7976]<=tmp[7875]*kernel[0]+tmp[7876]*kernel[1]+tmp[7877]*kernel[2]+tmp[7975]*kernel[3]+tmp[7976]*kernel[4]+tmp[7977]*kernel[5]+tmp[8075]*kernel[6]+tmp[8076]*kernel[7]+tmp[8077]*kernel[8];
				ans[7977]<=tmp[7876]*kernel[0]+tmp[7877]*kernel[1]+tmp[7878]*kernel[2]+tmp[7976]*kernel[3]+tmp[7977]*kernel[4]+tmp[7978]*kernel[5]+tmp[8076]*kernel[6]+tmp[8077]*kernel[7]+tmp[8078]*kernel[8];
				ans[7978]<=tmp[7877]*kernel[0]+tmp[7878]*kernel[1]+tmp[7879]*kernel[2]+tmp[7977]*kernel[3]+tmp[7978]*kernel[4]+tmp[7979]*kernel[5]+tmp[8077]*kernel[6]+tmp[8078]*kernel[7]+tmp[8079]*kernel[8];
				ans[7979]<=tmp[7878]*kernel[0]+tmp[7879]*kernel[1]+tmp[7880]*kernel[2]+tmp[7978]*kernel[3]+tmp[7979]*kernel[4]+tmp[7980]*kernel[5]+tmp[8078]*kernel[6]+tmp[8079]*kernel[7]+tmp[8080]*kernel[8];
				ans[7980]<=tmp[7879]*kernel[0]+tmp[7880]*kernel[1]+tmp[7881]*kernel[2]+tmp[7979]*kernel[3]+tmp[7980]*kernel[4]+tmp[7981]*kernel[5]+tmp[8079]*kernel[6]+tmp[8080]*kernel[7]+tmp[8081]*kernel[8];
				ans[7981]<=tmp[7880]*kernel[0]+tmp[7881]*kernel[1]+tmp[7882]*kernel[2]+tmp[7980]*kernel[3]+tmp[7981]*kernel[4]+tmp[7982]*kernel[5]+tmp[8080]*kernel[6]+tmp[8081]*kernel[7]+tmp[8082]*kernel[8];
				ans[7982]<=tmp[7881]*kernel[0]+tmp[7882]*kernel[1]+tmp[7883]*kernel[2]+tmp[7981]*kernel[3]+tmp[7982]*kernel[4]+tmp[7983]*kernel[5]+tmp[8081]*kernel[6]+tmp[8082]*kernel[7]+tmp[8083]*kernel[8];
				ans[7983]<=tmp[7882]*kernel[0]+tmp[7883]*kernel[1]+tmp[7884]*kernel[2]+tmp[7982]*kernel[3]+tmp[7983]*kernel[4]+tmp[7984]*kernel[5]+tmp[8082]*kernel[6]+tmp[8083]*kernel[7]+tmp[8084]*kernel[8];
				ans[7984]<=tmp[7883]*kernel[0]+tmp[7884]*kernel[1]+tmp[7885]*kernel[2]+tmp[7983]*kernel[3]+tmp[7984]*kernel[4]+tmp[7985]*kernel[5]+tmp[8083]*kernel[6]+tmp[8084]*kernel[7]+tmp[8085]*kernel[8];
				ans[7985]<=tmp[7884]*kernel[0]+tmp[7885]*kernel[1]+tmp[7886]*kernel[2]+tmp[7984]*kernel[3]+tmp[7985]*kernel[4]+tmp[7986]*kernel[5]+tmp[8084]*kernel[6]+tmp[8085]*kernel[7]+tmp[8086]*kernel[8];
				ans[7986]<=tmp[7885]*kernel[0]+tmp[7886]*kernel[1]+tmp[7887]*kernel[2]+tmp[7985]*kernel[3]+tmp[7986]*kernel[4]+tmp[7987]*kernel[5]+tmp[8085]*kernel[6]+tmp[8086]*kernel[7]+tmp[8087]*kernel[8];
				ans[7987]<=tmp[7886]*kernel[0]+tmp[7887]*kernel[1]+tmp[7888]*kernel[2]+tmp[7986]*kernel[3]+tmp[7987]*kernel[4]+tmp[7988]*kernel[5]+tmp[8086]*kernel[6]+tmp[8087]*kernel[7]+tmp[8088]*kernel[8];
				ans[7988]<=tmp[7887]*kernel[0]+tmp[7888]*kernel[1]+tmp[7889]*kernel[2]+tmp[7987]*kernel[3]+tmp[7988]*kernel[4]+tmp[7989]*kernel[5]+tmp[8087]*kernel[6]+tmp[8088]*kernel[7]+tmp[8089]*kernel[8];
				ans[7989]<=tmp[7888]*kernel[0]+tmp[7889]*kernel[1]+tmp[7890]*kernel[2]+tmp[7988]*kernel[3]+tmp[7989]*kernel[4]+tmp[7990]*kernel[5]+tmp[8088]*kernel[6]+tmp[8089]*kernel[7]+tmp[8090]*kernel[8];
				ans[7990]<=tmp[7889]*kernel[0]+tmp[7890]*kernel[1]+tmp[7891]*kernel[2]+tmp[7989]*kernel[3]+tmp[7990]*kernel[4]+tmp[7991]*kernel[5]+tmp[8089]*kernel[6]+tmp[8090]*kernel[7]+tmp[8091]*kernel[8];
				ans[7991]<=tmp[7890]*kernel[0]+tmp[7891]*kernel[1]+tmp[7892]*kernel[2]+tmp[7990]*kernel[3]+tmp[7991]*kernel[4]+tmp[7992]*kernel[5]+tmp[8090]*kernel[6]+tmp[8091]*kernel[7]+tmp[8092]*kernel[8];
				ans[7992]<=tmp[7891]*kernel[0]+tmp[7892]*kernel[1]+tmp[7893]*kernel[2]+tmp[7991]*kernel[3]+tmp[7992]*kernel[4]+tmp[7993]*kernel[5]+tmp[8091]*kernel[6]+tmp[8092]*kernel[7]+tmp[8093]*kernel[8];
				ans[7993]<=tmp[7892]*kernel[0]+tmp[7893]*kernel[1]+tmp[7894]*kernel[2]+tmp[7992]*kernel[3]+tmp[7993]*kernel[4]+tmp[7994]*kernel[5]+tmp[8092]*kernel[6]+tmp[8093]*kernel[7]+tmp[8094]*kernel[8];
				ans[7994]<=tmp[7893]*kernel[0]+tmp[7894]*kernel[1]+tmp[7895]*kernel[2]+tmp[7993]*kernel[3]+tmp[7994]*kernel[4]+tmp[7995]*kernel[5]+tmp[8093]*kernel[6]+tmp[8094]*kernel[7]+tmp[8095]*kernel[8];
				ans[7995]<=tmp[7894]*kernel[0]+tmp[7895]*kernel[1]+tmp[7896]*kernel[2]+tmp[7994]*kernel[3]+tmp[7995]*kernel[4]+tmp[7996]*kernel[5]+tmp[8094]*kernel[6]+tmp[8095]*kernel[7]+tmp[8096]*kernel[8];
				ans[7996]<=tmp[7895]*kernel[0]+tmp[7896]*kernel[1]+tmp[7897]*kernel[2]+tmp[7995]*kernel[3]+tmp[7996]*kernel[4]+tmp[7997]*kernel[5]+tmp[8095]*kernel[6]+tmp[8096]*kernel[7]+tmp[8097]*kernel[8];
				ans[7997]<=tmp[7896]*kernel[0]+tmp[7897]*kernel[1]+tmp[7898]*kernel[2]+tmp[7996]*kernel[3]+tmp[7997]*kernel[4]+tmp[7998]*kernel[5]+tmp[8096]*kernel[6]+tmp[8097]*kernel[7]+tmp[8098]*kernel[8];
				ans[7998]<=tmp[7897]*kernel[0]+tmp[7898]*kernel[1]+tmp[7899]*kernel[2]+tmp[7997]*kernel[3]+tmp[7998]*kernel[4]+tmp[7999]*kernel[5]+tmp[8097]*kernel[6]+tmp[8098]*kernel[7]+tmp[8099]*kernel[8];
				ans[7999]<=tmp[7898]*kernel[0]+tmp[7899]*kernel[1]+tmp[7998]*kernel[3]+tmp[7999]*kernel[4]+tmp[8098]*kernel[6]+tmp[8099]*kernel[7];
				ans[8000]<=tmp[7900]*kernel[1]+tmp[7901]*kernel[2]+tmp[8000]*kernel[4]+tmp[8001]*kernel[5]+tmp[8100]*kernel[7]+tmp[8101]*kernel[8];
				ans[8001]<=tmp[7900]*kernel[0]+tmp[7901]*kernel[1]+tmp[7902]*kernel[2]+tmp[8000]*kernel[3]+tmp[8001]*kernel[4]+tmp[8002]*kernel[5]+tmp[8100]*kernel[6]+tmp[8101]*kernel[7]+tmp[8102]*kernel[8];
				ans[8002]<=tmp[7901]*kernel[0]+tmp[7902]*kernel[1]+tmp[7903]*kernel[2]+tmp[8001]*kernel[3]+tmp[8002]*kernel[4]+tmp[8003]*kernel[5]+tmp[8101]*kernel[6]+tmp[8102]*kernel[7]+tmp[8103]*kernel[8];
				ans[8003]<=tmp[7902]*kernel[0]+tmp[7903]*kernel[1]+tmp[7904]*kernel[2]+tmp[8002]*kernel[3]+tmp[8003]*kernel[4]+tmp[8004]*kernel[5]+tmp[8102]*kernel[6]+tmp[8103]*kernel[7]+tmp[8104]*kernel[8];
				ans[8004]<=tmp[7903]*kernel[0]+tmp[7904]*kernel[1]+tmp[7905]*kernel[2]+tmp[8003]*kernel[3]+tmp[8004]*kernel[4]+tmp[8005]*kernel[5]+tmp[8103]*kernel[6]+tmp[8104]*kernel[7]+tmp[8105]*kernel[8];
				ans[8005]<=tmp[7904]*kernel[0]+tmp[7905]*kernel[1]+tmp[7906]*kernel[2]+tmp[8004]*kernel[3]+tmp[8005]*kernel[4]+tmp[8006]*kernel[5]+tmp[8104]*kernel[6]+tmp[8105]*kernel[7]+tmp[8106]*kernel[8];
				ans[8006]<=tmp[7905]*kernel[0]+tmp[7906]*kernel[1]+tmp[7907]*kernel[2]+tmp[8005]*kernel[3]+tmp[8006]*kernel[4]+tmp[8007]*kernel[5]+tmp[8105]*kernel[6]+tmp[8106]*kernel[7]+tmp[8107]*kernel[8];
				ans[8007]<=tmp[7906]*kernel[0]+tmp[7907]*kernel[1]+tmp[7908]*kernel[2]+tmp[8006]*kernel[3]+tmp[8007]*kernel[4]+tmp[8008]*kernel[5]+tmp[8106]*kernel[6]+tmp[8107]*kernel[7]+tmp[8108]*kernel[8];
				ans[8008]<=tmp[7907]*kernel[0]+tmp[7908]*kernel[1]+tmp[7909]*kernel[2]+tmp[8007]*kernel[3]+tmp[8008]*kernel[4]+tmp[8009]*kernel[5]+tmp[8107]*kernel[6]+tmp[8108]*kernel[7]+tmp[8109]*kernel[8];
				ans[8009]<=tmp[7908]*kernel[0]+tmp[7909]*kernel[1]+tmp[7910]*kernel[2]+tmp[8008]*kernel[3]+tmp[8009]*kernel[4]+tmp[8010]*kernel[5]+tmp[8108]*kernel[6]+tmp[8109]*kernel[7]+tmp[8110]*kernel[8];
				ans[8010]<=tmp[7909]*kernel[0]+tmp[7910]*kernel[1]+tmp[7911]*kernel[2]+tmp[8009]*kernel[3]+tmp[8010]*kernel[4]+tmp[8011]*kernel[5]+tmp[8109]*kernel[6]+tmp[8110]*kernel[7]+tmp[8111]*kernel[8];
				ans[8011]<=tmp[7910]*kernel[0]+tmp[7911]*kernel[1]+tmp[7912]*kernel[2]+tmp[8010]*kernel[3]+tmp[8011]*kernel[4]+tmp[8012]*kernel[5]+tmp[8110]*kernel[6]+tmp[8111]*kernel[7]+tmp[8112]*kernel[8];
				ans[8012]<=tmp[7911]*kernel[0]+tmp[7912]*kernel[1]+tmp[7913]*kernel[2]+tmp[8011]*kernel[3]+tmp[8012]*kernel[4]+tmp[8013]*kernel[5]+tmp[8111]*kernel[6]+tmp[8112]*kernel[7]+tmp[8113]*kernel[8];
				ans[8013]<=tmp[7912]*kernel[0]+tmp[7913]*kernel[1]+tmp[7914]*kernel[2]+tmp[8012]*kernel[3]+tmp[8013]*kernel[4]+tmp[8014]*kernel[5]+tmp[8112]*kernel[6]+tmp[8113]*kernel[7]+tmp[8114]*kernel[8];
				ans[8014]<=tmp[7913]*kernel[0]+tmp[7914]*kernel[1]+tmp[7915]*kernel[2]+tmp[8013]*kernel[3]+tmp[8014]*kernel[4]+tmp[8015]*kernel[5]+tmp[8113]*kernel[6]+tmp[8114]*kernel[7]+tmp[8115]*kernel[8];
				ans[8015]<=tmp[7914]*kernel[0]+tmp[7915]*kernel[1]+tmp[7916]*kernel[2]+tmp[8014]*kernel[3]+tmp[8015]*kernel[4]+tmp[8016]*kernel[5]+tmp[8114]*kernel[6]+tmp[8115]*kernel[7]+tmp[8116]*kernel[8];
				ans[8016]<=tmp[7915]*kernel[0]+tmp[7916]*kernel[1]+tmp[7917]*kernel[2]+tmp[8015]*kernel[3]+tmp[8016]*kernel[4]+tmp[8017]*kernel[5]+tmp[8115]*kernel[6]+tmp[8116]*kernel[7]+tmp[8117]*kernel[8];
				ans[8017]<=tmp[7916]*kernel[0]+tmp[7917]*kernel[1]+tmp[7918]*kernel[2]+tmp[8016]*kernel[3]+tmp[8017]*kernel[4]+tmp[8018]*kernel[5]+tmp[8116]*kernel[6]+tmp[8117]*kernel[7]+tmp[8118]*kernel[8];
				ans[8018]<=tmp[7917]*kernel[0]+tmp[7918]*kernel[1]+tmp[7919]*kernel[2]+tmp[8017]*kernel[3]+tmp[8018]*kernel[4]+tmp[8019]*kernel[5]+tmp[8117]*kernel[6]+tmp[8118]*kernel[7]+tmp[8119]*kernel[8];
				ans[8019]<=tmp[7918]*kernel[0]+tmp[7919]*kernel[1]+tmp[7920]*kernel[2]+tmp[8018]*kernel[3]+tmp[8019]*kernel[4]+tmp[8020]*kernel[5]+tmp[8118]*kernel[6]+tmp[8119]*kernel[7]+tmp[8120]*kernel[8];
				ans[8020]<=tmp[7919]*kernel[0]+tmp[7920]*kernel[1]+tmp[7921]*kernel[2]+tmp[8019]*kernel[3]+tmp[8020]*kernel[4]+tmp[8021]*kernel[5]+tmp[8119]*kernel[6]+tmp[8120]*kernel[7]+tmp[8121]*kernel[8];
				ans[8021]<=tmp[7920]*kernel[0]+tmp[7921]*kernel[1]+tmp[7922]*kernel[2]+tmp[8020]*kernel[3]+tmp[8021]*kernel[4]+tmp[8022]*kernel[5]+tmp[8120]*kernel[6]+tmp[8121]*kernel[7]+tmp[8122]*kernel[8];
				ans[8022]<=tmp[7921]*kernel[0]+tmp[7922]*kernel[1]+tmp[7923]*kernel[2]+tmp[8021]*kernel[3]+tmp[8022]*kernel[4]+tmp[8023]*kernel[5]+tmp[8121]*kernel[6]+tmp[8122]*kernel[7]+tmp[8123]*kernel[8];
				ans[8023]<=tmp[7922]*kernel[0]+tmp[7923]*kernel[1]+tmp[7924]*kernel[2]+tmp[8022]*kernel[3]+tmp[8023]*kernel[4]+tmp[8024]*kernel[5]+tmp[8122]*kernel[6]+tmp[8123]*kernel[7]+tmp[8124]*kernel[8];
				ans[8024]<=tmp[7923]*kernel[0]+tmp[7924]*kernel[1]+tmp[7925]*kernel[2]+tmp[8023]*kernel[3]+tmp[8024]*kernel[4]+tmp[8025]*kernel[5]+tmp[8123]*kernel[6]+tmp[8124]*kernel[7]+tmp[8125]*kernel[8];
				ans[8025]<=tmp[7924]*kernel[0]+tmp[7925]*kernel[1]+tmp[7926]*kernel[2]+tmp[8024]*kernel[3]+tmp[8025]*kernel[4]+tmp[8026]*kernel[5]+tmp[8124]*kernel[6]+tmp[8125]*kernel[7]+tmp[8126]*kernel[8];
				ans[8026]<=tmp[7925]*kernel[0]+tmp[7926]*kernel[1]+tmp[7927]*kernel[2]+tmp[8025]*kernel[3]+tmp[8026]*kernel[4]+tmp[8027]*kernel[5]+tmp[8125]*kernel[6]+tmp[8126]*kernel[7]+tmp[8127]*kernel[8];
				ans[8027]<=tmp[7926]*kernel[0]+tmp[7927]*kernel[1]+tmp[7928]*kernel[2]+tmp[8026]*kernel[3]+tmp[8027]*kernel[4]+tmp[8028]*kernel[5]+tmp[8126]*kernel[6]+tmp[8127]*kernel[7]+tmp[8128]*kernel[8];
				ans[8028]<=tmp[7927]*kernel[0]+tmp[7928]*kernel[1]+tmp[7929]*kernel[2]+tmp[8027]*kernel[3]+tmp[8028]*kernel[4]+tmp[8029]*kernel[5]+tmp[8127]*kernel[6]+tmp[8128]*kernel[7]+tmp[8129]*kernel[8];
				ans[8029]<=tmp[7928]*kernel[0]+tmp[7929]*kernel[1]+tmp[7930]*kernel[2]+tmp[8028]*kernel[3]+tmp[8029]*kernel[4]+tmp[8030]*kernel[5]+tmp[8128]*kernel[6]+tmp[8129]*kernel[7]+tmp[8130]*kernel[8];
				ans[8030]<=tmp[7929]*kernel[0]+tmp[7930]*kernel[1]+tmp[7931]*kernel[2]+tmp[8029]*kernel[3]+tmp[8030]*kernel[4]+tmp[8031]*kernel[5]+tmp[8129]*kernel[6]+tmp[8130]*kernel[7]+tmp[8131]*kernel[8];
				ans[8031]<=tmp[7930]*kernel[0]+tmp[7931]*kernel[1]+tmp[7932]*kernel[2]+tmp[8030]*kernel[3]+tmp[8031]*kernel[4]+tmp[8032]*kernel[5]+tmp[8130]*kernel[6]+tmp[8131]*kernel[7]+tmp[8132]*kernel[8];
				ans[8032]<=tmp[7931]*kernel[0]+tmp[7932]*kernel[1]+tmp[7933]*kernel[2]+tmp[8031]*kernel[3]+tmp[8032]*kernel[4]+tmp[8033]*kernel[5]+tmp[8131]*kernel[6]+tmp[8132]*kernel[7]+tmp[8133]*kernel[8];
				ans[8033]<=tmp[7932]*kernel[0]+tmp[7933]*kernel[1]+tmp[7934]*kernel[2]+tmp[8032]*kernel[3]+tmp[8033]*kernel[4]+tmp[8034]*kernel[5]+tmp[8132]*kernel[6]+tmp[8133]*kernel[7]+tmp[8134]*kernel[8];
				ans[8034]<=tmp[7933]*kernel[0]+tmp[7934]*kernel[1]+tmp[7935]*kernel[2]+tmp[8033]*kernel[3]+tmp[8034]*kernel[4]+tmp[8035]*kernel[5]+tmp[8133]*kernel[6]+tmp[8134]*kernel[7]+tmp[8135]*kernel[8];
				ans[8035]<=tmp[7934]*kernel[0]+tmp[7935]*kernel[1]+tmp[7936]*kernel[2]+tmp[8034]*kernel[3]+tmp[8035]*kernel[4]+tmp[8036]*kernel[5]+tmp[8134]*kernel[6]+tmp[8135]*kernel[7]+tmp[8136]*kernel[8];
				ans[8036]<=tmp[7935]*kernel[0]+tmp[7936]*kernel[1]+tmp[7937]*kernel[2]+tmp[8035]*kernel[3]+tmp[8036]*kernel[4]+tmp[8037]*kernel[5]+tmp[8135]*kernel[6]+tmp[8136]*kernel[7]+tmp[8137]*kernel[8];
				ans[8037]<=tmp[7936]*kernel[0]+tmp[7937]*kernel[1]+tmp[7938]*kernel[2]+tmp[8036]*kernel[3]+tmp[8037]*kernel[4]+tmp[8038]*kernel[5]+tmp[8136]*kernel[6]+tmp[8137]*kernel[7]+tmp[8138]*kernel[8];
				ans[8038]<=tmp[7937]*kernel[0]+tmp[7938]*kernel[1]+tmp[7939]*kernel[2]+tmp[8037]*kernel[3]+tmp[8038]*kernel[4]+tmp[8039]*kernel[5]+tmp[8137]*kernel[6]+tmp[8138]*kernel[7]+tmp[8139]*kernel[8];
				ans[8039]<=tmp[7938]*kernel[0]+tmp[7939]*kernel[1]+tmp[7940]*kernel[2]+tmp[8038]*kernel[3]+tmp[8039]*kernel[4]+tmp[8040]*kernel[5]+tmp[8138]*kernel[6]+tmp[8139]*kernel[7]+tmp[8140]*kernel[8];
				ans[8040]<=tmp[7939]*kernel[0]+tmp[7940]*kernel[1]+tmp[7941]*kernel[2]+tmp[8039]*kernel[3]+tmp[8040]*kernel[4]+tmp[8041]*kernel[5]+tmp[8139]*kernel[6]+tmp[8140]*kernel[7]+tmp[8141]*kernel[8];
				ans[8041]<=tmp[7940]*kernel[0]+tmp[7941]*kernel[1]+tmp[7942]*kernel[2]+tmp[8040]*kernel[3]+tmp[8041]*kernel[4]+tmp[8042]*kernel[5]+tmp[8140]*kernel[6]+tmp[8141]*kernel[7]+tmp[8142]*kernel[8];
				ans[8042]<=tmp[7941]*kernel[0]+tmp[7942]*kernel[1]+tmp[7943]*kernel[2]+tmp[8041]*kernel[3]+tmp[8042]*kernel[4]+tmp[8043]*kernel[5]+tmp[8141]*kernel[6]+tmp[8142]*kernel[7]+tmp[8143]*kernel[8];
				ans[8043]<=tmp[7942]*kernel[0]+tmp[7943]*kernel[1]+tmp[7944]*kernel[2]+tmp[8042]*kernel[3]+tmp[8043]*kernel[4]+tmp[8044]*kernel[5]+tmp[8142]*kernel[6]+tmp[8143]*kernel[7]+tmp[8144]*kernel[8];
				ans[8044]<=tmp[7943]*kernel[0]+tmp[7944]*kernel[1]+tmp[7945]*kernel[2]+tmp[8043]*kernel[3]+tmp[8044]*kernel[4]+tmp[8045]*kernel[5]+tmp[8143]*kernel[6]+tmp[8144]*kernel[7]+tmp[8145]*kernel[8];
				ans[8045]<=tmp[7944]*kernel[0]+tmp[7945]*kernel[1]+tmp[7946]*kernel[2]+tmp[8044]*kernel[3]+tmp[8045]*kernel[4]+tmp[8046]*kernel[5]+tmp[8144]*kernel[6]+tmp[8145]*kernel[7]+tmp[8146]*kernel[8];
				ans[8046]<=tmp[7945]*kernel[0]+tmp[7946]*kernel[1]+tmp[7947]*kernel[2]+tmp[8045]*kernel[3]+tmp[8046]*kernel[4]+tmp[8047]*kernel[5]+tmp[8145]*kernel[6]+tmp[8146]*kernel[7]+tmp[8147]*kernel[8];
				ans[8047]<=tmp[7946]*kernel[0]+tmp[7947]*kernel[1]+tmp[7948]*kernel[2]+tmp[8046]*kernel[3]+tmp[8047]*kernel[4]+tmp[8048]*kernel[5]+tmp[8146]*kernel[6]+tmp[8147]*kernel[7]+tmp[8148]*kernel[8];
				ans[8048]<=tmp[7947]*kernel[0]+tmp[7948]*kernel[1]+tmp[7949]*kernel[2]+tmp[8047]*kernel[3]+tmp[8048]*kernel[4]+tmp[8049]*kernel[5]+tmp[8147]*kernel[6]+tmp[8148]*kernel[7]+tmp[8149]*kernel[8];
				ans[8049]<=tmp[7948]*kernel[0]+tmp[7949]*kernel[1]+tmp[7950]*kernel[2]+tmp[8048]*kernel[3]+tmp[8049]*kernel[4]+tmp[8050]*kernel[5]+tmp[8148]*kernel[6]+tmp[8149]*kernel[7]+tmp[8150]*kernel[8];
				ans[8050]<=tmp[7949]*kernel[0]+tmp[7950]*kernel[1]+tmp[7951]*kernel[2]+tmp[8049]*kernel[3]+tmp[8050]*kernel[4]+tmp[8051]*kernel[5]+tmp[8149]*kernel[6]+tmp[8150]*kernel[7]+tmp[8151]*kernel[8];
				ans[8051]<=tmp[7950]*kernel[0]+tmp[7951]*kernel[1]+tmp[7952]*kernel[2]+tmp[8050]*kernel[3]+tmp[8051]*kernel[4]+tmp[8052]*kernel[5]+tmp[8150]*kernel[6]+tmp[8151]*kernel[7]+tmp[8152]*kernel[8];
				ans[8052]<=tmp[7951]*kernel[0]+tmp[7952]*kernel[1]+tmp[7953]*kernel[2]+tmp[8051]*kernel[3]+tmp[8052]*kernel[4]+tmp[8053]*kernel[5]+tmp[8151]*kernel[6]+tmp[8152]*kernel[7]+tmp[8153]*kernel[8];
				ans[8053]<=tmp[7952]*kernel[0]+tmp[7953]*kernel[1]+tmp[7954]*kernel[2]+tmp[8052]*kernel[3]+tmp[8053]*kernel[4]+tmp[8054]*kernel[5]+tmp[8152]*kernel[6]+tmp[8153]*kernel[7]+tmp[8154]*kernel[8];
				ans[8054]<=tmp[7953]*kernel[0]+tmp[7954]*kernel[1]+tmp[7955]*kernel[2]+tmp[8053]*kernel[3]+tmp[8054]*kernel[4]+tmp[8055]*kernel[5]+tmp[8153]*kernel[6]+tmp[8154]*kernel[7]+tmp[8155]*kernel[8];
				ans[8055]<=tmp[7954]*kernel[0]+tmp[7955]*kernel[1]+tmp[7956]*kernel[2]+tmp[8054]*kernel[3]+tmp[8055]*kernel[4]+tmp[8056]*kernel[5]+tmp[8154]*kernel[6]+tmp[8155]*kernel[7]+tmp[8156]*kernel[8];
				ans[8056]<=tmp[7955]*kernel[0]+tmp[7956]*kernel[1]+tmp[7957]*kernel[2]+tmp[8055]*kernel[3]+tmp[8056]*kernel[4]+tmp[8057]*kernel[5]+tmp[8155]*kernel[6]+tmp[8156]*kernel[7]+tmp[8157]*kernel[8];
				ans[8057]<=tmp[7956]*kernel[0]+tmp[7957]*kernel[1]+tmp[7958]*kernel[2]+tmp[8056]*kernel[3]+tmp[8057]*kernel[4]+tmp[8058]*kernel[5]+tmp[8156]*kernel[6]+tmp[8157]*kernel[7]+tmp[8158]*kernel[8];
				ans[8058]<=tmp[7957]*kernel[0]+tmp[7958]*kernel[1]+tmp[7959]*kernel[2]+tmp[8057]*kernel[3]+tmp[8058]*kernel[4]+tmp[8059]*kernel[5]+tmp[8157]*kernel[6]+tmp[8158]*kernel[7]+tmp[8159]*kernel[8];
				ans[8059]<=tmp[7958]*kernel[0]+tmp[7959]*kernel[1]+tmp[7960]*kernel[2]+tmp[8058]*kernel[3]+tmp[8059]*kernel[4]+tmp[8060]*kernel[5]+tmp[8158]*kernel[6]+tmp[8159]*kernel[7]+tmp[8160]*kernel[8];
				ans[8060]<=tmp[7959]*kernel[0]+tmp[7960]*kernel[1]+tmp[7961]*kernel[2]+tmp[8059]*kernel[3]+tmp[8060]*kernel[4]+tmp[8061]*kernel[5]+tmp[8159]*kernel[6]+tmp[8160]*kernel[7]+tmp[8161]*kernel[8];
				ans[8061]<=tmp[7960]*kernel[0]+tmp[7961]*kernel[1]+tmp[7962]*kernel[2]+tmp[8060]*kernel[3]+tmp[8061]*kernel[4]+tmp[8062]*kernel[5]+tmp[8160]*kernel[6]+tmp[8161]*kernel[7]+tmp[8162]*kernel[8];
				ans[8062]<=tmp[7961]*kernel[0]+tmp[7962]*kernel[1]+tmp[7963]*kernel[2]+tmp[8061]*kernel[3]+tmp[8062]*kernel[4]+tmp[8063]*kernel[5]+tmp[8161]*kernel[6]+tmp[8162]*kernel[7]+tmp[8163]*kernel[8];
				ans[8063]<=tmp[7962]*kernel[0]+tmp[7963]*kernel[1]+tmp[7964]*kernel[2]+tmp[8062]*kernel[3]+tmp[8063]*kernel[4]+tmp[8064]*kernel[5]+tmp[8162]*kernel[6]+tmp[8163]*kernel[7]+tmp[8164]*kernel[8];
				ans[8064]<=tmp[7963]*kernel[0]+tmp[7964]*kernel[1]+tmp[7965]*kernel[2]+tmp[8063]*kernel[3]+tmp[8064]*kernel[4]+tmp[8065]*kernel[5]+tmp[8163]*kernel[6]+tmp[8164]*kernel[7]+tmp[8165]*kernel[8];
				ans[8065]<=tmp[7964]*kernel[0]+tmp[7965]*kernel[1]+tmp[7966]*kernel[2]+tmp[8064]*kernel[3]+tmp[8065]*kernel[4]+tmp[8066]*kernel[5]+tmp[8164]*kernel[6]+tmp[8165]*kernel[7]+tmp[8166]*kernel[8];
				ans[8066]<=tmp[7965]*kernel[0]+tmp[7966]*kernel[1]+tmp[7967]*kernel[2]+tmp[8065]*kernel[3]+tmp[8066]*kernel[4]+tmp[8067]*kernel[5]+tmp[8165]*kernel[6]+tmp[8166]*kernel[7]+tmp[8167]*kernel[8];
				ans[8067]<=tmp[7966]*kernel[0]+tmp[7967]*kernel[1]+tmp[7968]*kernel[2]+tmp[8066]*kernel[3]+tmp[8067]*kernel[4]+tmp[8068]*kernel[5]+tmp[8166]*kernel[6]+tmp[8167]*kernel[7]+tmp[8168]*kernel[8];
				ans[8068]<=tmp[7967]*kernel[0]+tmp[7968]*kernel[1]+tmp[7969]*kernel[2]+tmp[8067]*kernel[3]+tmp[8068]*kernel[4]+tmp[8069]*kernel[5]+tmp[8167]*kernel[6]+tmp[8168]*kernel[7]+tmp[8169]*kernel[8];
				ans[8069]<=tmp[7968]*kernel[0]+tmp[7969]*kernel[1]+tmp[7970]*kernel[2]+tmp[8068]*kernel[3]+tmp[8069]*kernel[4]+tmp[8070]*kernel[5]+tmp[8168]*kernel[6]+tmp[8169]*kernel[7]+tmp[8170]*kernel[8];
				ans[8070]<=tmp[7969]*kernel[0]+tmp[7970]*kernel[1]+tmp[7971]*kernel[2]+tmp[8069]*kernel[3]+tmp[8070]*kernel[4]+tmp[8071]*kernel[5]+tmp[8169]*kernel[6]+tmp[8170]*kernel[7]+tmp[8171]*kernel[8];
				ans[8071]<=tmp[7970]*kernel[0]+tmp[7971]*kernel[1]+tmp[7972]*kernel[2]+tmp[8070]*kernel[3]+tmp[8071]*kernel[4]+tmp[8072]*kernel[5]+tmp[8170]*kernel[6]+tmp[8171]*kernel[7]+tmp[8172]*kernel[8];
				ans[8072]<=tmp[7971]*kernel[0]+tmp[7972]*kernel[1]+tmp[7973]*kernel[2]+tmp[8071]*kernel[3]+tmp[8072]*kernel[4]+tmp[8073]*kernel[5]+tmp[8171]*kernel[6]+tmp[8172]*kernel[7]+tmp[8173]*kernel[8];
				ans[8073]<=tmp[7972]*kernel[0]+tmp[7973]*kernel[1]+tmp[7974]*kernel[2]+tmp[8072]*kernel[3]+tmp[8073]*kernel[4]+tmp[8074]*kernel[5]+tmp[8172]*kernel[6]+tmp[8173]*kernel[7]+tmp[8174]*kernel[8];
				ans[8074]<=tmp[7973]*kernel[0]+tmp[7974]*kernel[1]+tmp[7975]*kernel[2]+tmp[8073]*kernel[3]+tmp[8074]*kernel[4]+tmp[8075]*kernel[5]+tmp[8173]*kernel[6]+tmp[8174]*kernel[7]+tmp[8175]*kernel[8];
				ans[8075]<=tmp[7974]*kernel[0]+tmp[7975]*kernel[1]+tmp[7976]*kernel[2]+tmp[8074]*kernel[3]+tmp[8075]*kernel[4]+tmp[8076]*kernel[5]+tmp[8174]*kernel[6]+tmp[8175]*kernel[7]+tmp[8176]*kernel[8];
				ans[8076]<=tmp[7975]*kernel[0]+tmp[7976]*kernel[1]+tmp[7977]*kernel[2]+tmp[8075]*kernel[3]+tmp[8076]*kernel[4]+tmp[8077]*kernel[5]+tmp[8175]*kernel[6]+tmp[8176]*kernel[7]+tmp[8177]*kernel[8];
				ans[8077]<=tmp[7976]*kernel[0]+tmp[7977]*kernel[1]+tmp[7978]*kernel[2]+tmp[8076]*kernel[3]+tmp[8077]*kernel[4]+tmp[8078]*kernel[5]+tmp[8176]*kernel[6]+tmp[8177]*kernel[7]+tmp[8178]*kernel[8];
				ans[8078]<=tmp[7977]*kernel[0]+tmp[7978]*kernel[1]+tmp[7979]*kernel[2]+tmp[8077]*kernel[3]+tmp[8078]*kernel[4]+tmp[8079]*kernel[5]+tmp[8177]*kernel[6]+tmp[8178]*kernel[7]+tmp[8179]*kernel[8];
				ans[8079]<=tmp[7978]*kernel[0]+tmp[7979]*kernel[1]+tmp[7980]*kernel[2]+tmp[8078]*kernel[3]+tmp[8079]*kernel[4]+tmp[8080]*kernel[5]+tmp[8178]*kernel[6]+tmp[8179]*kernel[7]+tmp[8180]*kernel[8];
				ans[8080]<=tmp[7979]*kernel[0]+tmp[7980]*kernel[1]+tmp[7981]*kernel[2]+tmp[8079]*kernel[3]+tmp[8080]*kernel[4]+tmp[8081]*kernel[5]+tmp[8179]*kernel[6]+tmp[8180]*kernel[7]+tmp[8181]*kernel[8];
				ans[8081]<=tmp[7980]*kernel[0]+tmp[7981]*kernel[1]+tmp[7982]*kernel[2]+tmp[8080]*kernel[3]+tmp[8081]*kernel[4]+tmp[8082]*kernel[5]+tmp[8180]*kernel[6]+tmp[8181]*kernel[7]+tmp[8182]*kernel[8];
				ans[8082]<=tmp[7981]*kernel[0]+tmp[7982]*kernel[1]+tmp[7983]*kernel[2]+tmp[8081]*kernel[3]+tmp[8082]*kernel[4]+tmp[8083]*kernel[5]+tmp[8181]*kernel[6]+tmp[8182]*kernel[7]+tmp[8183]*kernel[8];
				ans[8083]<=tmp[7982]*kernel[0]+tmp[7983]*kernel[1]+tmp[7984]*kernel[2]+tmp[8082]*kernel[3]+tmp[8083]*kernel[4]+tmp[8084]*kernel[5]+tmp[8182]*kernel[6]+tmp[8183]*kernel[7]+tmp[8184]*kernel[8];
				ans[8084]<=tmp[7983]*kernel[0]+tmp[7984]*kernel[1]+tmp[7985]*kernel[2]+tmp[8083]*kernel[3]+tmp[8084]*kernel[4]+tmp[8085]*kernel[5]+tmp[8183]*kernel[6]+tmp[8184]*kernel[7]+tmp[8185]*kernel[8];
				ans[8085]<=tmp[7984]*kernel[0]+tmp[7985]*kernel[1]+tmp[7986]*kernel[2]+tmp[8084]*kernel[3]+tmp[8085]*kernel[4]+tmp[8086]*kernel[5]+tmp[8184]*kernel[6]+tmp[8185]*kernel[7]+tmp[8186]*kernel[8];
				ans[8086]<=tmp[7985]*kernel[0]+tmp[7986]*kernel[1]+tmp[7987]*kernel[2]+tmp[8085]*kernel[3]+tmp[8086]*kernel[4]+tmp[8087]*kernel[5]+tmp[8185]*kernel[6]+tmp[8186]*kernel[7]+tmp[8187]*kernel[8];
				ans[8087]<=tmp[7986]*kernel[0]+tmp[7987]*kernel[1]+tmp[7988]*kernel[2]+tmp[8086]*kernel[3]+tmp[8087]*kernel[4]+tmp[8088]*kernel[5]+tmp[8186]*kernel[6]+tmp[8187]*kernel[7]+tmp[8188]*kernel[8];
				ans[8088]<=tmp[7987]*kernel[0]+tmp[7988]*kernel[1]+tmp[7989]*kernel[2]+tmp[8087]*kernel[3]+tmp[8088]*kernel[4]+tmp[8089]*kernel[5]+tmp[8187]*kernel[6]+tmp[8188]*kernel[7]+tmp[8189]*kernel[8];
				ans[8089]<=tmp[7988]*kernel[0]+tmp[7989]*kernel[1]+tmp[7990]*kernel[2]+tmp[8088]*kernel[3]+tmp[8089]*kernel[4]+tmp[8090]*kernel[5]+tmp[8188]*kernel[6]+tmp[8189]*kernel[7]+tmp[8190]*kernel[8];
				ans[8090]<=tmp[7989]*kernel[0]+tmp[7990]*kernel[1]+tmp[7991]*kernel[2]+tmp[8089]*kernel[3]+tmp[8090]*kernel[4]+tmp[8091]*kernel[5]+tmp[8189]*kernel[6]+tmp[8190]*kernel[7]+tmp[8191]*kernel[8];
				ans[8091]<=tmp[7990]*kernel[0]+tmp[7991]*kernel[1]+tmp[7992]*kernel[2]+tmp[8090]*kernel[3]+tmp[8091]*kernel[4]+tmp[8092]*kernel[5]+tmp[8190]*kernel[6]+tmp[8191]*kernel[7]+tmp[8192]*kernel[8];
				ans[8092]<=tmp[7991]*kernel[0]+tmp[7992]*kernel[1]+tmp[7993]*kernel[2]+tmp[8091]*kernel[3]+tmp[8092]*kernel[4]+tmp[8093]*kernel[5]+tmp[8191]*kernel[6]+tmp[8192]*kernel[7]+tmp[8193]*kernel[8];
				ans[8093]<=tmp[7992]*kernel[0]+tmp[7993]*kernel[1]+tmp[7994]*kernel[2]+tmp[8092]*kernel[3]+tmp[8093]*kernel[4]+tmp[8094]*kernel[5]+tmp[8192]*kernel[6]+tmp[8193]*kernel[7]+tmp[8194]*kernel[8];
				ans[8094]<=tmp[7993]*kernel[0]+tmp[7994]*kernel[1]+tmp[7995]*kernel[2]+tmp[8093]*kernel[3]+tmp[8094]*kernel[4]+tmp[8095]*kernel[5]+tmp[8193]*kernel[6]+tmp[8194]*kernel[7]+tmp[8195]*kernel[8];
				ans[8095]<=tmp[7994]*kernel[0]+tmp[7995]*kernel[1]+tmp[7996]*kernel[2]+tmp[8094]*kernel[3]+tmp[8095]*kernel[4]+tmp[8096]*kernel[5]+tmp[8194]*kernel[6]+tmp[8195]*kernel[7]+tmp[8196]*kernel[8];
				ans[8096]<=tmp[7995]*kernel[0]+tmp[7996]*kernel[1]+tmp[7997]*kernel[2]+tmp[8095]*kernel[3]+tmp[8096]*kernel[4]+tmp[8097]*kernel[5]+tmp[8195]*kernel[6]+tmp[8196]*kernel[7]+tmp[8197]*kernel[8];
				ans[8097]<=tmp[7996]*kernel[0]+tmp[7997]*kernel[1]+tmp[7998]*kernel[2]+tmp[8096]*kernel[3]+tmp[8097]*kernel[4]+tmp[8098]*kernel[5]+tmp[8196]*kernel[6]+tmp[8197]*kernel[7]+tmp[8198]*kernel[8];
				ans[8098]<=tmp[7997]*kernel[0]+tmp[7998]*kernel[1]+tmp[7999]*kernel[2]+tmp[8097]*kernel[3]+tmp[8098]*kernel[4]+tmp[8099]*kernel[5]+tmp[8197]*kernel[6]+tmp[8198]*kernel[7]+tmp[8199]*kernel[8];
				ans[8099]<=tmp[7998]*kernel[0]+tmp[7999]*kernel[1]+tmp[8098]*kernel[3]+tmp[8099]*kernel[4]+tmp[8198]*kernel[6]+tmp[8199]*kernel[7];
				ans[8100]<=tmp[8000]*kernel[1]+tmp[8001]*kernel[2]+tmp[8100]*kernel[4]+tmp[8101]*kernel[5]+tmp[8200]*kernel[7]+tmp[8201]*kernel[8];
				ans[8101]<=tmp[8000]*kernel[0]+tmp[8001]*kernel[1]+tmp[8002]*kernel[2]+tmp[8100]*kernel[3]+tmp[8101]*kernel[4]+tmp[8102]*kernel[5]+tmp[8200]*kernel[6]+tmp[8201]*kernel[7]+tmp[8202]*kernel[8];
				ans[8102]<=tmp[8001]*kernel[0]+tmp[8002]*kernel[1]+tmp[8003]*kernel[2]+tmp[8101]*kernel[3]+tmp[8102]*kernel[4]+tmp[8103]*kernel[5]+tmp[8201]*kernel[6]+tmp[8202]*kernel[7]+tmp[8203]*kernel[8];
				ans[8103]<=tmp[8002]*kernel[0]+tmp[8003]*kernel[1]+tmp[8004]*kernel[2]+tmp[8102]*kernel[3]+tmp[8103]*kernel[4]+tmp[8104]*kernel[5]+tmp[8202]*kernel[6]+tmp[8203]*kernel[7]+tmp[8204]*kernel[8];
				ans[8104]<=tmp[8003]*kernel[0]+tmp[8004]*kernel[1]+tmp[8005]*kernel[2]+tmp[8103]*kernel[3]+tmp[8104]*kernel[4]+tmp[8105]*kernel[5]+tmp[8203]*kernel[6]+tmp[8204]*kernel[7]+tmp[8205]*kernel[8];
				ans[8105]<=tmp[8004]*kernel[0]+tmp[8005]*kernel[1]+tmp[8006]*kernel[2]+tmp[8104]*kernel[3]+tmp[8105]*kernel[4]+tmp[8106]*kernel[5]+tmp[8204]*kernel[6]+tmp[8205]*kernel[7]+tmp[8206]*kernel[8];
				ans[8106]<=tmp[8005]*kernel[0]+tmp[8006]*kernel[1]+tmp[8007]*kernel[2]+tmp[8105]*kernel[3]+tmp[8106]*kernel[4]+tmp[8107]*kernel[5]+tmp[8205]*kernel[6]+tmp[8206]*kernel[7]+tmp[8207]*kernel[8];
				ans[8107]<=tmp[8006]*kernel[0]+tmp[8007]*kernel[1]+tmp[8008]*kernel[2]+tmp[8106]*kernel[3]+tmp[8107]*kernel[4]+tmp[8108]*kernel[5]+tmp[8206]*kernel[6]+tmp[8207]*kernel[7]+tmp[8208]*kernel[8];
				ans[8108]<=tmp[8007]*kernel[0]+tmp[8008]*kernel[1]+tmp[8009]*kernel[2]+tmp[8107]*kernel[3]+tmp[8108]*kernel[4]+tmp[8109]*kernel[5]+tmp[8207]*kernel[6]+tmp[8208]*kernel[7]+tmp[8209]*kernel[8];
				ans[8109]<=tmp[8008]*kernel[0]+tmp[8009]*kernel[1]+tmp[8010]*kernel[2]+tmp[8108]*kernel[3]+tmp[8109]*kernel[4]+tmp[8110]*kernel[5]+tmp[8208]*kernel[6]+tmp[8209]*kernel[7]+tmp[8210]*kernel[8];
				ans[8110]<=tmp[8009]*kernel[0]+tmp[8010]*kernel[1]+tmp[8011]*kernel[2]+tmp[8109]*kernel[3]+tmp[8110]*kernel[4]+tmp[8111]*kernel[5]+tmp[8209]*kernel[6]+tmp[8210]*kernel[7]+tmp[8211]*kernel[8];
				ans[8111]<=tmp[8010]*kernel[0]+tmp[8011]*kernel[1]+tmp[8012]*kernel[2]+tmp[8110]*kernel[3]+tmp[8111]*kernel[4]+tmp[8112]*kernel[5]+tmp[8210]*kernel[6]+tmp[8211]*kernel[7]+tmp[8212]*kernel[8];
				ans[8112]<=tmp[8011]*kernel[0]+tmp[8012]*kernel[1]+tmp[8013]*kernel[2]+tmp[8111]*kernel[3]+tmp[8112]*kernel[4]+tmp[8113]*kernel[5]+tmp[8211]*kernel[6]+tmp[8212]*kernel[7]+tmp[8213]*kernel[8];
				ans[8113]<=tmp[8012]*kernel[0]+tmp[8013]*kernel[1]+tmp[8014]*kernel[2]+tmp[8112]*kernel[3]+tmp[8113]*kernel[4]+tmp[8114]*kernel[5]+tmp[8212]*kernel[6]+tmp[8213]*kernel[7]+tmp[8214]*kernel[8];
				ans[8114]<=tmp[8013]*kernel[0]+tmp[8014]*kernel[1]+tmp[8015]*kernel[2]+tmp[8113]*kernel[3]+tmp[8114]*kernel[4]+tmp[8115]*kernel[5]+tmp[8213]*kernel[6]+tmp[8214]*kernel[7]+tmp[8215]*kernel[8];
				ans[8115]<=tmp[8014]*kernel[0]+tmp[8015]*kernel[1]+tmp[8016]*kernel[2]+tmp[8114]*kernel[3]+tmp[8115]*kernel[4]+tmp[8116]*kernel[5]+tmp[8214]*kernel[6]+tmp[8215]*kernel[7]+tmp[8216]*kernel[8];
				ans[8116]<=tmp[8015]*kernel[0]+tmp[8016]*kernel[1]+tmp[8017]*kernel[2]+tmp[8115]*kernel[3]+tmp[8116]*kernel[4]+tmp[8117]*kernel[5]+tmp[8215]*kernel[6]+tmp[8216]*kernel[7]+tmp[8217]*kernel[8];
				ans[8117]<=tmp[8016]*kernel[0]+tmp[8017]*kernel[1]+tmp[8018]*kernel[2]+tmp[8116]*kernel[3]+tmp[8117]*kernel[4]+tmp[8118]*kernel[5]+tmp[8216]*kernel[6]+tmp[8217]*kernel[7]+tmp[8218]*kernel[8];
				ans[8118]<=tmp[8017]*kernel[0]+tmp[8018]*kernel[1]+tmp[8019]*kernel[2]+tmp[8117]*kernel[3]+tmp[8118]*kernel[4]+tmp[8119]*kernel[5]+tmp[8217]*kernel[6]+tmp[8218]*kernel[7]+tmp[8219]*kernel[8];
				ans[8119]<=tmp[8018]*kernel[0]+tmp[8019]*kernel[1]+tmp[8020]*kernel[2]+tmp[8118]*kernel[3]+tmp[8119]*kernel[4]+tmp[8120]*kernel[5]+tmp[8218]*kernel[6]+tmp[8219]*kernel[7]+tmp[8220]*kernel[8];
				ans[8120]<=tmp[8019]*kernel[0]+tmp[8020]*kernel[1]+tmp[8021]*kernel[2]+tmp[8119]*kernel[3]+tmp[8120]*kernel[4]+tmp[8121]*kernel[5]+tmp[8219]*kernel[6]+tmp[8220]*kernel[7]+tmp[8221]*kernel[8];
				ans[8121]<=tmp[8020]*kernel[0]+tmp[8021]*kernel[1]+tmp[8022]*kernel[2]+tmp[8120]*kernel[3]+tmp[8121]*kernel[4]+tmp[8122]*kernel[5]+tmp[8220]*kernel[6]+tmp[8221]*kernel[7]+tmp[8222]*kernel[8];
				ans[8122]<=tmp[8021]*kernel[0]+tmp[8022]*kernel[1]+tmp[8023]*kernel[2]+tmp[8121]*kernel[3]+tmp[8122]*kernel[4]+tmp[8123]*kernel[5]+tmp[8221]*kernel[6]+tmp[8222]*kernel[7]+tmp[8223]*kernel[8];
				ans[8123]<=tmp[8022]*kernel[0]+tmp[8023]*kernel[1]+tmp[8024]*kernel[2]+tmp[8122]*kernel[3]+tmp[8123]*kernel[4]+tmp[8124]*kernel[5]+tmp[8222]*kernel[6]+tmp[8223]*kernel[7]+tmp[8224]*kernel[8];
				ans[8124]<=tmp[8023]*kernel[0]+tmp[8024]*kernel[1]+tmp[8025]*kernel[2]+tmp[8123]*kernel[3]+tmp[8124]*kernel[4]+tmp[8125]*kernel[5]+tmp[8223]*kernel[6]+tmp[8224]*kernel[7]+tmp[8225]*kernel[8];
				ans[8125]<=tmp[8024]*kernel[0]+tmp[8025]*kernel[1]+tmp[8026]*kernel[2]+tmp[8124]*kernel[3]+tmp[8125]*kernel[4]+tmp[8126]*kernel[5]+tmp[8224]*kernel[6]+tmp[8225]*kernel[7]+tmp[8226]*kernel[8];
				ans[8126]<=tmp[8025]*kernel[0]+tmp[8026]*kernel[1]+tmp[8027]*kernel[2]+tmp[8125]*kernel[3]+tmp[8126]*kernel[4]+tmp[8127]*kernel[5]+tmp[8225]*kernel[6]+tmp[8226]*kernel[7]+tmp[8227]*kernel[8];
				ans[8127]<=tmp[8026]*kernel[0]+tmp[8027]*kernel[1]+tmp[8028]*kernel[2]+tmp[8126]*kernel[3]+tmp[8127]*kernel[4]+tmp[8128]*kernel[5]+tmp[8226]*kernel[6]+tmp[8227]*kernel[7]+tmp[8228]*kernel[8];
				ans[8128]<=tmp[8027]*kernel[0]+tmp[8028]*kernel[1]+tmp[8029]*kernel[2]+tmp[8127]*kernel[3]+tmp[8128]*kernel[4]+tmp[8129]*kernel[5]+tmp[8227]*kernel[6]+tmp[8228]*kernel[7]+tmp[8229]*kernel[8];
				ans[8129]<=tmp[8028]*kernel[0]+tmp[8029]*kernel[1]+tmp[8030]*kernel[2]+tmp[8128]*kernel[3]+tmp[8129]*kernel[4]+tmp[8130]*kernel[5]+tmp[8228]*kernel[6]+tmp[8229]*kernel[7]+tmp[8230]*kernel[8];
				ans[8130]<=tmp[8029]*kernel[0]+tmp[8030]*kernel[1]+tmp[8031]*kernel[2]+tmp[8129]*kernel[3]+tmp[8130]*kernel[4]+tmp[8131]*kernel[5]+tmp[8229]*kernel[6]+tmp[8230]*kernel[7]+tmp[8231]*kernel[8];
				ans[8131]<=tmp[8030]*kernel[0]+tmp[8031]*kernel[1]+tmp[8032]*kernel[2]+tmp[8130]*kernel[3]+tmp[8131]*kernel[4]+tmp[8132]*kernel[5]+tmp[8230]*kernel[6]+tmp[8231]*kernel[7]+tmp[8232]*kernel[8];
				ans[8132]<=tmp[8031]*kernel[0]+tmp[8032]*kernel[1]+tmp[8033]*kernel[2]+tmp[8131]*kernel[3]+tmp[8132]*kernel[4]+tmp[8133]*kernel[5]+tmp[8231]*kernel[6]+tmp[8232]*kernel[7]+tmp[8233]*kernel[8];
				ans[8133]<=tmp[8032]*kernel[0]+tmp[8033]*kernel[1]+tmp[8034]*kernel[2]+tmp[8132]*kernel[3]+tmp[8133]*kernel[4]+tmp[8134]*kernel[5]+tmp[8232]*kernel[6]+tmp[8233]*kernel[7]+tmp[8234]*kernel[8];
				ans[8134]<=tmp[8033]*kernel[0]+tmp[8034]*kernel[1]+tmp[8035]*kernel[2]+tmp[8133]*kernel[3]+tmp[8134]*kernel[4]+tmp[8135]*kernel[5]+tmp[8233]*kernel[6]+tmp[8234]*kernel[7]+tmp[8235]*kernel[8];
				ans[8135]<=tmp[8034]*kernel[0]+tmp[8035]*kernel[1]+tmp[8036]*kernel[2]+tmp[8134]*kernel[3]+tmp[8135]*kernel[4]+tmp[8136]*kernel[5]+tmp[8234]*kernel[6]+tmp[8235]*kernel[7]+tmp[8236]*kernel[8];
				ans[8136]<=tmp[8035]*kernel[0]+tmp[8036]*kernel[1]+tmp[8037]*kernel[2]+tmp[8135]*kernel[3]+tmp[8136]*kernel[4]+tmp[8137]*kernel[5]+tmp[8235]*kernel[6]+tmp[8236]*kernel[7]+tmp[8237]*kernel[8];
				ans[8137]<=tmp[8036]*kernel[0]+tmp[8037]*kernel[1]+tmp[8038]*kernel[2]+tmp[8136]*kernel[3]+tmp[8137]*kernel[4]+tmp[8138]*kernel[5]+tmp[8236]*kernel[6]+tmp[8237]*kernel[7]+tmp[8238]*kernel[8];
				ans[8138]<=tmp[8037]*kernel[0]+tmp[8038]*kernel[1]+tmp[8039]*kernel[2]+tmp[8137]*kernel[3]+tmp[8138]*kernel[4]+tmp[8139]*kernel[5]+tmp[8237]*kernel[6]+tmp[8238]*kernel[7]+tmp[8239]*kernel[8];
				ans[8139]<=tmp[8038]*kernel[0]+tmp[8039]*kernel[1]+tmp[8040]*kernel[2]+tmp[8138]*kernel[3]+tmp[8139]*kernel[4]+tmp[8140]*kernel[5]+tmp[8238]*kernel[6]+tmp[8239]*kernel[7]+tmp[8240]*kernel[8];
				ans[8140]<=tmp[8039]*kernel[0]+tmp[8040]*kernel[1]+tmp[8041]*kernel[2]+tmp[8139]*kernel[3]+tmp[8140]*kernel[4]+tmp[8141]*kernel[5]+tmp[8239]*kernel[6]+tmp[8240]*kernel[7]+tmp[8241]*kernel[8];
				ans[8141]<=tmp[8040]*kernel[0]+tmp[8041]*kernel[1]+tmp[8042]*kernel[2]+tmp[8140]*kernel[3]+tmp[8141]*kernel[4]+tmp[8142]*kernel[5]+tmp[8240]*kernel[6]+tmp[8241]*kernel[7]+tmp[8242]*kernel[8];
				ans[8142]<=tmp[8041]*kernel[0]+tmp[8042]*kernel[1]+tmp[8043]*kernel[2]+tmp[8141]*kernel[3]+tmp[8142]*kernel[4]+tmp[8143]*kernel[5]+tmp[8241]*kernel[6]+tmp[8242]*kernel[7]+tmp[8243]*kernel[8];
				ans[8143]<=tmp[8042]*kernel[0]+tmp[8043]*kernel[1]+tmp[8044]*kernel[2]+tmp[8142]*kernel[3]+tmp[8143]*kernel[4]+tmp[8144]*kernel[5]+tmp[8242]*kernel[6]+tmp[8243]*kernel[7]+tmp[8244]*kernel[8];
				ans[8144]<=tmp[8043]*kernel[0]+tmp[8044]*kernel[1]+tmp[8045]*kernel[2]+tmp[8143]*kernel[3]+tmp[8144]*kernel[4]+tmp[8145]*kernel[5]+tmp[8243]*kernel[6]+tmp[8244]*kernel[7]+tmp[8245]*kernel[8];
				ans[8145]<=tmp[8044]*kernel[0]+tmp[8045]*kernel[1]+tmp[8046]*kernel[2]+tmp[8144]*kernel[3]+tmp[8145]*kernel[4]+tmp[8146]*kernel[5]+tmp[8244]*kernel[6]+tmp[8245]*kernel[7]+tmp[8246]*kernel[8];
				ans[8146]<=tmp[8045]*kernel[0]+tmp[8046]*kernel[1]+tmp[8047]*kernel[2]+tmp[8145]*kernel[3]+tmp[8146]*kernel[4]+tmp[8147]*kernel[5]+tmp[8245]*kernel[6]+tmp[8246]*kernel[7]+tmp[8247]*kernel[8];
				ans[8147]<=tmp[8046]*kernel[0]+tmp[8047]*kernel[1]+tmp[8048]*kernel[2]+tmp[8146]*kernel[3]+tmp[8147]*kernel[4]+tmp[8148]*kernel[5]+tmp[8246]*kernel[6]+tmp[8247]*kernel[7]+tmp[8248]*kernel[8];
				ans[8148]<=tmp[8047]*kernel[0]+tmp[8048]*kernel[1]+tmp[8049]*kernel[2]+tmp[8147]*kernel[3]+tmp[8148]*kernel[4]+tmp[8149]*kernel[5]+tmp[8247]*kernel[6]+tmp[8248]*kernel[7]+tmp[8249]*kernel[8];
				ans[8149]<=tmp[8048]*kernel[0]+tmp[8049]*kernel[1]+tmp[8050]*kernel[2]+tmp[8148]*kernel[3]+tmp[8149]*kernel[4]+tmp[8150]*kernel[5]+tmp[8248]*kernel[6]+tmp[8249]*kernel[7]+tmp[8250]*kernel[8];
				ans[8150]<=tmp[8049]*kernel[0]+tmp[8050]*kernel[1]+tmp[8051]*kernel[2]+tmp[8149]*kernel[3]+tmp[8150]*kernel[4]+tmp[8151]*kernel[5]+tmp[8249]*kernel[6]+tmp[8250]*kernel[7]+tmp[8251]*kernel[8];
				ans[8151]<=tmp[8050]*kernel[0]+tmp[8051]*kernel[1]+tmp[8052]*kernel[2]+tmp[8150]*kernel[3]+tmp[8151]*kernel[4]+tmp[8152]*kernel[5]+tmp[8250]*kernel[6]+tmp[8251]*kernel[7]+tmp[8252]*kernel[8];
				ans[8152]<=tmp[8051]*kernel[0]+tmp[8052]*kernel[1]+tmp[8053]*kernel[2]+tmp[8151]*kernel[3]+tmp[8152]*kernel[4]+tmp[8153]*kernel[5]+tmp[8251]*kernel[6]+tmp[8252]*kernel[7]+tmp[8253]*kernel[8];
				ans[8153]<=tmp[8052]*kernel[0]+tmp[8053]*kernel[1]+tmp[8054]*kernel[2]+tmp[8152]*kernel[3]+tmp[8153]*kernel[4]+tmp[8154]*kernel[5]+tmp[8252]*kernel[6]+tmp[8253]*kernel[7]+tmp[8254]*kernel[8];
				ans[8154]<=tmp[8053]*kernel[0]+tmp[8054]*kernel[1]+tmp[8055]*kernel[2]+tmp[8153]*kernel[3]+tmp[8154]*kernel[4]+tmp[8155]*kernel[5]+tmp[8253]*kernel[6]+tmp[8254]*kernel[7]+tmp[8255]*kernel[8];
				ans[8155]<=tmp[8054]*kernel[0]+tmp[8055]*kernel[1]+tmp[8056]*kernel[2]+tmp[8154]*kernel[3]+tmp[8155]*kernel[4]+tmp[8156]*kernel[5]+tmp[8254]*kernel[6]+tmp[8255]*kernel[7]+tmp[8256]*kernel[8];
				ans[8156]<=tmp[8055]*kernel[0]+tmp[8056]*kernel[1]+tmp[8057]*kernel[2]+tmp[8155]*kernel[3]+tmp[8156]*kernel[4]+tmp[8157]*kernel[5]+tmp[8255]*kernel[6]+tmp[8256]*kernel[7]+tmp[8257]*kernel[8];
				ans[8157]<=tmp[8056]*kernel[0]+tmp[8057]*kernel[1]+tmp[8058]*kernel[2]+tmp[8156]*kernel[3]+tmp[8157]*kernel[4]+tmp[8158]*kernel[5]+tmp[8256]*kernel[6]+tmp[8257]*kernel[7]+tmp[8258]*kernel[8];
				ans[8158]<=tmp[8057]*kernel[0]+tmp[8058]*kernel[1]+tmp[8059]*kernel[2]+tmp[8157]*kernel[3]+tmp[8158]*kernel[4]+tmp[8159]*kernel[5]+tmp[8257]*kernel[6]+tmp[8258]*kernel[7]+tmp[8259]*kernel[8];
				ans[8159]<=tmp[8058]*kernel[0]+tmp[8059]*kernel[1]+tmp[8060]*kernel[2]+tmp[8158]*kernel[3]+tmp[8159]*kernel[4]+tmp[8160]*kernel[5]+tmp[8258]*kernel[6]+tmp[8259]*kernel[7]+tmp[8260]*kernel[8];
				ans[8160]<=tmp[8059]*kernel[0]+tmp[8060]*kernel[1]+tmp[8061]*kernel[2]+tmp[8159]*kernel[3]+tmp[8160]*kernel[4]+tmp[8161]*kernel[5]+tmp[8259]*kernel[6]+tmp[8260]*kernel[7]+tmp[8261]*kernel[8];
				ans[8161]<=tmp[8060]*kernel[0]+tmp[8061]*kernel[1]+tmp[8062]*kernel[2]+tmp[8160]*kernel[3]+tmp[8161]*kernel[4]+tmp[8162]*kernel[5]+tmp[8260]*kernel[6]+tmp[8261]*kernel[7]+tmp[8262]*kernel[8];
				ans[8162]<=tmp[8061]*kernel[0]+tmp[8062]*kernel[1]+tmp[8063]*kernel[2]+tmp[8161]*kernel[3]+tmp[8162]*kernel[4]+tmp[8163]*kernel[5]+tmp[8261]*kernel[6]+tmp[8262]*kernel[7]+tmp[8263]*kernel[8];
				ans[8163]<=tmp[8062]*kernel[0]+tmp[8063]*kernel[1]+tmp[8064]*kernel[2]+tmp[8162]*kernel[3]+tmp[8163]*kernel[4]+tmp[8164]*kernel[5]+tmp[8262]*kernel[6]+tmp[8263]*kernel[7]+tmp[8264]*kernel[8];
				ans[8164]<=tmp[8063]*kernel[0]+tmp[8064]*kernel[1]+tmp[8065]*kernel[2]+tmp[8163]*kernel[3]+tmp[8164]*kernel[4]+tmp[8165]*kernel[5]+tmp[8263]*kernel[6]+tmp[8264]*kernel[7]+tmp[8265]*kernel[8];
				ans[8165]<=tmp[8064]*kernel[0]+tmp[8065]*kernel[1]+tmp[8066]*kernel[2]+tmp[8164]*kernel[3]+tmp[8165]*kernel[4]+tmp[8166]*kernel[5]+tmp[8264]*kernel[6]+tmp[8265]*kernel[7]+tmp[8266]*kernel[8];
				ans[8166]<=tmp[8065]*kernel[0]+tmp[8066]*kernel[1]+tmp[8067]*kernel[2]+tmp[8165]*kernel[3]+tmp[8166]*kernel[4]+tmp[8167]*kernel[5]+tmp[8265]*kernel[6]+tmp[8266]*kernel[7]+tmp[8267]*kernel[8];
				ans[8167]<=tmp[8066]*kernel[0]+tmp[8067]*kernel[1]+tmp[8068]*kernel[2]+tmp[8166]*kernel[3]+tmp[8167]*kernel[4]+tmp[8168]*kernel[5]+tmp[8266]*kernel[6]+tmp[8267]*kernel[7]+tmp[8268]*kernel[8];
				ans[8168]<=tmp[8067]*kernel[0]+tmp[8068]*kernel[1]+tmp[8069]*kernel[2]+tmp[8167]*kernel[3]+tmp[8168]*kernel[4]+tmp[8169]*kernel[5]+tmp[8267]*kernel[6]+tmp[8268]*kernel[7]+tmp[8269]*kernel[8];
				ans[8169]<=tmp[8068]*kernel[0]+tmp[8069]*kernel[1]+tmp[8070]*kernel[2]+tmp[8168]*kernel[3]+tmp[8169]*kernel[4]+tmp[8170]*kernel[5]+tmp[8268]*kernel[6]+tmp[8269]*kernel[7]+tmp[8270]*kernel[8];
				ans[8170]<=tmp[8069]*kernel[0]+tmp[8070]*kernel[1]+tmp[8071]*kernel[2]+tmp[8169]*kernel[3]+tmp[8170]*kernel[4]+tmp[8171]*kernel[5]+tmp[8269]*kernel[6]+tmp[8270]*kernel[7]+tmp[8271]*kernel[8];
				ans[8171]<=tmp[8070]*kernel[0]+tmp[8071]*kernel[1]+tmp[8072]*kernel[2]+tmp[8170]*kernel[3]+tmp[8171]*kernel[4]+tmp[8172]*kernel[5]+tmp[8270]*kernel[6]+tmp[8271]*kernel[7]+tmp[8272]*kernel[8];
				ans[8172]<=tmp[8071]*kernel[0]+tmp[8072]*kernel[1]+tmp[8073]*kernel[2]+tmp[8171]*kernel[3]+tmp[8172]*kernel[4]+tmp[8173]*kernel[5]+tmp[8271]*kernel[6]+tmp[8272]*kernel[7]+tmp[8273]*kernel[8];
				ans[8173]<=tmp[8072]*kernel[0]+tmp[8073]*kernel[1]+tmp[8074]*kernel[2]+tmp[8172]*kernel[3]+tmp[8173]*kernel[4]+tmp[8174]*kernel[5]+tmp[8272]*kernel[6]+tmp[8273]*kernel[7]+tmp[8274]*kernel[8];
				ans[8174]<=tmp[8073]*kernel[0]+tmp[8074]*kernel[1]+tmp[8075]*kernel[2]+tmp[8173]*kernel[3]+tmp[8174]*kernel[4]+tmp[8175]*kernel[5]+tmp[8273]*kernel[6]+tmp[8274]*kernel[7]+tmp[8275]*kernel[8];
				ans[8175]<=tmp[8074]*kernel[0]+tmp[8075]*kernel[1]+tmp[8076]*kernel[2]+tmp[8174]*kernel[3]+tmp[8175]*kernel[4]+tmp[8176]*kernel[5]+tmp[8274]*kernel[6]+tmp[8275]*kernel[7]+tmp[8276]*kernel[8];
				ans[8176]<=tmp[8075]*kernel[0]+tmp[8076]*kernel[1]+tmp[8077]*kernel[2]+tmp[8175]*kernel[3]+tmp[8176]*kernel[4]+tmp[8177]*kernel[5]+tmp[8275]*kernel[6]+tmp[8276]*kernel[7]+tmp[8277]*kernel[8];
				ans[8177]<=tmp[8076]*kernel[0]+tmp[8077]*kernel[1]+tmp[8078]*kernel[2]+tmp[8176]*kernel[3]+tmp[8177]*kernel[4]+tmp[8178]*kernel[5]+tmp[8276]*kernel[6]+tmp[8277]*kernel[7]+tmp[8278]*kernel[8];
				ans[8178]<=tmp[8077]*kernel[0]+tmp[8078]*kernel[1]+tmp[8079]*kernel[2]+tmp[8177]*kernel[3]+tmp[8178]*kernel[4]+tmp[8179]*kernel[5]+tmp[8277]*kernel[6]+tmp[8278]*kernel[7]+tmp[8279]*kernel[8];
				ans[8179]<=tmp[8078]*kernel[0]+tmp[8079]*kernel[1]+tmp[8080]*kernel[2]+tmp[8178]*kernel[3]+tmp[8179]*kernel[4]+tmp[8180]*kernel[5]+tmp[8278]*kernel[6]+tmp[8279]*kernel[7]+tmp[8280]*kernel[8];
				ans[8180]<=tmp[8079]*kernel[0]+tmp[8080]*kernel[1]+tmp[8081]*kernel[2]+tmp[8179]*kernel[3]+tmp[8180]*kernel[4]+tmp[8181]*kernel[5]+tmp[8279]*kernel[6]+tmp[8280]*kernel[7]+tmp[8281]*kernel[8];
				ans[8181]<=tmp[8080]*kernel[0]+tmp[8081]*kernel[1]+tmp[8082]*kernel[2]+tmp[8180]*kernel[3]+tmp[8181]*kernel[4]+tmp[8182]*kernel[5]+tmp[8280]*kernel[6]+tmp[8281]*kernel[7]+tmp[8282]*kernel[8];
				ans[8182]<=tmp[8081]*kernel[0]+tmp[8082]*kernel[1]+tmp[8083]*kernel[2]+tmp[8181]*kernel[3]+tmp[8182]*kernel[4]+tmp[8183]*kernel[5]+tmp[8281]*kernel[6]+tmp[8282]*kernel[7]+tmp[8283]*kernel[8];
				ans[8183]<=tmp[8082]*kernel[0]+tmp[8083]*kernel[1]+tmp[8084]*kernel[2]+tmp[8182]*kernel[3]+tmp[8183]*kernel[4]+tmp[8184]*kernel[5]+tmp[8282]*kernel[6]+tmp[8283]*kernel[7]+tmp[8284]*kernel[8];
				ans[8184]<=tmp[8083]*kernel[0]+tmp[8084]*kernel[1]+tmp[8085]*kernel[2]+tmp[8183]*kernel[3]+tmp[8184]*kernel[4]+tmp[8185]*kernel[5]+tmp[8283]*kernel[6]+tmp[8284]*kernel[7]+tmp[8285]*kernel[8];
				ans[8185]<=tmp[8084]*kernel[0]+tmp[8085]*kernel[1]+tmp[8086]*kernel[2]+tmp[8184]*kernel[3]+tmp[8185]*kernel[4]+tmp[8186]*kernel[5]+tmp[8284]*kernel[6]+tmp[8285]*kernel[7]+tmp[8286]*kernel[8];
				ans[8186]<=tmp[8085]*kernel[0]+tmp[8086]*kernel[1]+tmp[8087]*kernel[2]+tmp[8185]*kernel[3]+tmp[8186]*kernel[4]+tmp[8187]*kernel[5]+tmp[8285]*kernel[6]+tmp[8286]*kernel[7]+tmp[8287]*kernel[8];
				ans[8187]<=tmp[8086]*kernel[0]+tmp[8087]*kernel[1]+tmp[8088]*kernel[2]+tmp[8186]*kernel[3]+tmp[8187]*kernel[4]+tmp[8188]*kernel[5]+tmp[8286]*kernel[6]+tmp[8287]*kernel[7]+tmp[8288]*kernel[8];
				ans[8188]<=tmp[8087]*kernel[0]+tmp[8088]*kernel[1]+tmp[8089]*kernel[2]+tmp[8187]*kernel[3]+tmp[8188]*kernel[4]+tmp[8189]*kernel[5]+tmp[8287]*kernel[6]+tmp[8288]*kernel[7]+tmp[8289]*kernel[8];
				ans[8189]<=tmp[8088]*kernel[0]+tmp[8089]*kernel[1]+tmp[8090]*kernel[2]+tmp[8188]*kernel[3]+tmp[8189]*kernel[4]+tmp[8190]*kernel[5]+tmp[8288]*kernel[6]+tmp[8289]*kernel[7]+tmp[8290]*kernel[8];
				ans[8190]<=tmp[8089]*kernel[0]+tmp[8090]*kernel[1]+tmp[8091]*kernel[2]+tmp[8189]*kernel[3]+tmp[8190]*kernel[4]+tmp[8191]*kernel[5]+tmp[8289]*kernel[6]+tmp[8290]*kernel[7]+tmp[8291]*kernel[8];
				ans[8191]<=tmp[8090]*kernel[0]+tmp[8091]*kernel[1]+tmp[8092]*kernel[2]+tmp[8190]*kernel[3]+tmp[8191]*kernel[4]+tmp[8192]*kernel[5]+tmp[8290]*kernel[6]+tmp[8291]*kernel[7]+tmp[8292]*kernel[8];
				ans[8192]<=tmp[8091]*kernel[0]+tmp[8092]*kernel[1]+tmp[8093]*kernel[2]+tmp[8191]*kernel[3]+tmp[8192]*kernel[4]+tmp[8193]*kernel[5]+tmp[8291]*kernel[6]+tmp[8292]*kernel[7]+tmp[8293]*kernel[8];
				ans[8193]<=tmp[8092]*kernel[0]+tmp[8093]*kernel[1]+tmp[8094]*kernel[2]+tmp[8192]*kernel[3]+tmp[8193]*kernel[4]+tmp[8194]*kernel[5]+tmp[8292]*kernel[6]+tmp[8293]*kernel[7]+tmp[8294]*kernel[8];
				ans[8194]<=tmp[8093]*kernel[0]+tmp[8094]*kernel[1]+tmp[8095]*kernel[2]+tmp[8193]*kernel[3]+tmp[8194]*kernel[4]+tmp[8195]*kernel[5]+tmp[8293]*kernel[6]+tmp[8294]*kernel[7]+tmp[8295]*kernel[8];
				ans[8195]<=tmp[8094]*kernel[0]+tmp[8095]*kernel[1]+tmp[8096]*kernel[2]+tmp[8194]*kernel[3]+tmp[8195]*kernel[4]+tmp[8196]*kernel[5]+tmp[8294]*kernel[6]+tmp[8295]*kernel[7]+tmp[8296]*kernel[8];
				ans[8196]<=tmp[8095]*kernel[0]+tmp[8096]*kernel[1]+tmp[8097]*kernel[2]+tmp[8195]*kernel[3]+tmp[8196]*kernel[4]+tmp[8197]*kernel[5]+tmp[8295]*kernel[6]+tmp[8296]*kernel[7]+tmp[8297]*kernel[8];
				ans[8197]<=tmp[8096]*kernel[0]+tmp[8097]*kernel[1]+tmp[8098]*kernel[2]+tmp[8196]*kernel[3]+tmp[8197]*kernel[4]+tmp[8198]*kernel[5]+tmp[8296]*kernel[6]+tmp[8297]*kernel[7]+tmp[8298]*kernel[8];
				ans[8198]<=tmp[8097]*kernel[0]+tmp[8098]*kernel[1]+tmp[8099]*kernel[2]+tmp[8197]*kernel[3]+tmp[8198]*kernel[4]+tmp[8199]*kernel[5]+tmp[8297]*kernel[6]+tmp[8298]*kernel[7]+tmp[8299]*kernel[8];
				ans[8199]<=tmp[8098]*kernel[0]+tmp[8099]*kernel[1]+tmp[8198]*kernel[3]+tmp[8199]*kernel[4]+tmp[8298]*kernel[6]+tmp[8299]*kernel[7];
				ans[8200]<=tmp[8100]*kernel[1]+tmp[8101]*kernel[2]+tmp[8200]*kernel[4]+tmp[8201]*kernel[5]+tmp[8300]*kernel[7]+tmp[8301]*kernel[8];
				ans[8201]<=tmp[8100]*kernel[0]+tmp[8101]*kernel[1]+tmp[8102]*kernel[2]+tmp[8200]*kernel[3]+tmp[8201]*kernel[4]+tmp[8202]*kernel[5]+tmp[8300]*kernel[6]+tmp[8301]*kernel[7]+tmp[8302]*kernel[8];
				ans[8202]<=tmp[8101]*kernel[0]+tmp[8102]*kernel[1]+tmp[8103]*kernel[2]+tmp[8201]*kernel[3]+tmp[8202]*kernel[4]+tmp[8203]*kernel[5]+tmp[8301]*kernel[6]+tmp[8302]*kernel[7]+tmp[8303]*kernel[8];
				ans[8203]<=tmp[8102]*kernel[0]+tmp[8103]*kernel[1]+tmp[8104]*kernel[2]+tmp[8202]*kernel[3]+tmp[8203]*kernel[4]+tmp[8204]*kernel[5]+tmp[8302]*kernel[6]+tmp[8303]*kernel[7]+tmp[8304]*kernel[8];
				ans[8204]<=tmp[8103]*kernel[0]+tmp[8104]*kernel[1]+tmp[8105]*kernel[2]+tmp[8203]*kernel[3]+tmp[8204]*kernel[4]+tmp[8205]*kernel[5]+tmp[8303]*kernel[6]+tmp[8304]*kernel[7]+tmp[8305]*kernel[8];
				ans[8205]<=tmp[8104]*kernel[0]+tmp[8105]*kernel[1]+tmp[8106]*kernel[2]+tmp[8204]*kernel[3]+tmp[8205]*kernel[4]+tmp[8206]*kernel[5]+tmp[8304]*kernel[6]+tmp[8305]*kernel[7]+tmp[8306]*kernel[8];
				ans[8206]<=tmp[8105]*kernel[0]+tmp[8106]*kernel[1]+tmp[8107]*kernel[2]+tmp[8205]*kernel[3]+tmp[8206]*kernel[4]+tmp[8207]*kernel[5]+tmp[8305]*kernel[6]+tmp[8306]*kernel[7]+tmp[8307]*kernel[8];
				ans[8207]<=tmp[8106]*kernel[0]+tmp[8107]*kernel[1]+tmp[8108]*kernel[2]+tmp[8206]*kernel[3]+tmp[8207]*kernel[4]+tmp[8208]*kernel[5]+tmp[8306]*kernel[6]+tmp[8307]*kernel[7]+tmp[8308]*kernel[8];
				ans[8208]<=tmp[8107]*kernel[0]+tmp[8108]*kernel[1]+tmp[8109]*kernel[2]+tmp[8207]*kernel[3]+tmp[8208]*kernel[4]+tmp[8209]*kernel[5]+tmp[8307]*kernel[6]+tmp[8308]*kernel[7]+tmp[8309]*kernel[8];
				ans[8209]<=tmp[8108]*kernel[0]+tmp[8109]*kernel[1]+tmp[8110]*kernel[2]+tmp[8208]*kernel[3]+tmp[8209]*kernel[4]+tmp[8210]*kernel[5]+tmp[8308]*kernel[6]+tmp[8309]*kernel[7]+tmp[8310]*kernel[8];
				ans[8210]<=tmp[8109]*kernel[0]+tmp[8110]*kernel[1]+tmp[8111]*kernel[2]+tmp[8209]*kernel[3]+tmp[8210]*kernel[4]+tmp[8211]*kernel[5]+tmp[8309]*kernel[6]+tmp[8310]*kernel[7]+tmp[8311]*kernel[8];
				ans[8211]<=tmp[8110]*kernel[0]+tmp[8111]*kernel[1]+tmp[8112]*kernel[2]+tmp[8210]*kernel[3]+tmp[8211]*kernel[4]+tmp[8212]*kernel[5]+tmp[8310]*kernel[6]+tmp[8311]*kernel[7]+tmp[8312]*kernel[8];
				ans[8212]<=tmp[8111]*kernel[0]+tmp[8112]*kernel[1]+tmp[8113]*kernel[2]+tmp[8211]*kernel[3]+tmp[8212]*kernel[4]+tmp[8213]*kernel[5]+tmp[8311]*kernel[6]+tmp[8312]*kernel[7]+tmp[8313]*kernel[8];
				ans[8213]<=tmp[8112]*kernel[0]+tmp[8113]*kernel[1]+tmp[8114]*kernel[2]+tmp[8212]*kernel[3]+tmp[8213]*kernel[4]+tmp[8214]*kernel[5]+tmp[8312]*kernel[6]+tmp[8313]*kernel[7]+tmp[8314]*kernel[8];
				ans[8214]<=tmp[8113]*kernel[0]+tmp[8114]*kernel[1]+tmp[8115]*kernel[2]+tmp[8213]*kernel[3]+tmp[8214]*kernel[4]+tmp[8215]*kernel[5]+tmp[8313]*kernel[6]+tmp[8314]*kernel[7]+tmp[8315]*kernel[8];
				ans[8215]<=tmp[8114]*kernel[0]+tmp[8115]*kernel[1]+tmp[8116]*kernel[2]+tmp[8214]*kernel[3]+tmp[8215]*kernel[4]+tmp[8216]*kernel[5]+tmp[8314]*kernel[6]+tmp[8315]*kernel[7]+tmp[8316]*kernel[8];
				ans[8216]<=tmp[8115]*kernel[0]+tmp[8116]*kernel[1]+tmp[8117]*kernel[2]+tmp[8215]*kernel[3]+tmp[8216]*kernel[4]+tmp[8217]*kernel[5]+tmp[8315]*kernel[6]+tmp[8316]*kernel[7]+tmp[8317]*kernel[8];
				ans[8217]<=tmp[8116]*kernel[0]+tmp[8117]*kernel[1]+tmp[8118]*kernel[2]+tmp[8216]*kernel[3]+tmp[8217]*kernel[4]+tmp[8218]*kernel[5]+tmp[8316]*kernel[6]+tmp[8317]*kernel[7]+tmp[8318]*kernel[8];
				ans[8218]<=tmp[8117]*kernel[0]+tmp[8118]*kernel[1]+tmp[8119]*kernel[2]+tmp[8217]*kernel[3]+tmp[8218]*kernel[4]+tmp[8219]*kernel[5]+tmp[8317]*kernel[6]+tmp[8318]*kernel[7]+tmp[8319]*kernel[8];
				ans[8219]<=tmp[8118]*kernel[0]+tmp[8119]*kernel[1]+tmp[8120]*kernel[2]+tmp[8218]*kernel[3]+tmp[8219]*kernel[4]+tmp[8220]*kernel[5]+tmp[8318]*kernel[6]+tmp[8319]*kernel[7]+tmp[8320]*kernel[8];
				ans[8220]<=tmp[8119]*kernel[0]+tmp[8120]*kernel[1]+tmp[8121]*kernel[2]+tmp[8219]*kernel[3]+tmp[8220]*kernel[4]+tmp[8221]*kernel[5]+tmp[8319]*kernel[6]+tmp[8320]*kernel[7]+tmp[8321]*kernel[8];
				ans[8221]<=tmp[8120]*kernel[0]+tmp[8121]*kernel[1]+tmp[8122]*kernel[2]+tmp[8220]*kernel[3]+tmp[8221]*kernel[4]+tmp[8222]*kernel[5]+tmp[8320]*kernel[6]+tmp[8321]*kernel[7]+tmp[8322]*kernel[8];
				ans[8222]<=tmp[8121]*kernel[0]+tmp[8122]*kernel[1]+tmp[8123]*kernel[2]+tmp[8221]*kernel[3]+tmp[8222]*kernel[4]+tmp[8223]*kernel[5]+tmp[8321]*kernel[6]+tmp[8322]*kernel[7]+tmp[8323]*kernel[8];
				ans[8223]<=tmp[8122]*kernel[0]+tmp[8123]*kernel[1]+tmp[8124]*kernel[2]+tmp[8222]*kernel[3]+tmp[8223]*kernel[4]+tmp[8224]*kernel[5]+tmp[8322]*kernel[6]+tmp[8323]*kernel[7]+tmp[8324]*kernel[8];
				ans[8224]<=tmp[8123]*kernel[0]+tmp[8124]*kernel[1]+tmp[8125]*kernel[2]+tmp[8223]*kernel[3]+tmp[8224]*kernel[4]+tmp[8225]*kernel[5]+tmp[8323]*kernel[6]+tmp[8324]*kernel[7]+tmp[8325]*kernel[8];
				ans[8225]<=tmp[8124]*kernel[0]+tmp[8125]*kernel[1]+tmp[8126]*kernel[2]+tmp[8224]*kernel[3]+tmp[8225]*kernel[4]+tmp[8226]*kernel[5]+tmp[8324]*kernel[6]+tmp[8325]*kernel[7]+tmp[8326]*kernel[8];
				ans[8226]<=tmp[8125]*kernel[0]+tmp[8126]*kernel[1]+tmp[8127]*kernel[2]+tmp[8225]*kernel[3]+tmp[8226]*kernel[4]+tmp[8227]*kernel[5]+tmp[8325]*kernel[6]+tmp[8326]*kernel[7]+tmp[8327]*kernel[8];
				ans[8227]<=tmp[8126]*kernel[0]+tmp[8127]*kernel[1]+tmp[8128]*kernel[2]+tmp[8226]*kernel[3]+tmp[8227]*kernel[4]+tmp[8228]*kernel[5]+tmp[8326]*kernel[6]+tmp[8327]*kernel[7]+tmp[8328]*kernel[8];
				ans[8228]<=tmp[8127]*kernel[0]+tmp[8128]*kernel[1]+tmp[8129]*kernel[2]+tmp[8227]*kernel[3]+tmp[8228]*kernel[4]+tmp[8229]*kernel[5]+tmp[8327]*kernel[6]+tmp[8328]*kernel[7]+tmp[8329]*kernel[8];
				ans[8229]<=tmp[8128]*kernel[0]+tmp[8129]*kernel[1]+tmp[8130]*kernel[2]+tmp[8228]*kernel[3]+tmp[8229]*kernel[4]+tmp[8230]*kernel[5]+tmp[8328]*kernel[6]+tmp[8329]*kernel[7]+tmp[8330]*kernel[8];
				ans[8230]<=tmp[8129]*kernel[0]+tmp[8130]*kernel[1]+tmp[8131]*kernel[2]+tmp[8229]*kernel[3]+tmp[8230]*kernel[4]+tmp[8231]*kernel[5]+tmp[8329]*kernel[6]+tmp[8330]*kernel[7]+tmp[8331]*kernel[8];
				ans[8231]<=tmp[8130]*kernel[0]+tmp[8131]*kernel[1]+tmp[8132]*kernel[2]+tmp[8230]*kernel[3]+tmp[8231]*kernel[4]+tmp[8232]*kernel[5]+tmp[8330]*kernel[6]+tmp[8331]*kernel[7]+tmp[8332]*kernel[8];
				ans[8232]<=tmp[8131]*kernel[0]+tmp[8132]*kernel[1]+tmp[8133]*kernel[2]+tmp[8231]*kernel[3]+tmp[8232]*kernel[4]+tmp[8233]*kernel[5]+tmp[8331]*kernel[6]+tmp[8332]*kernel[7]+tmp[8333]*kernel[8];
				ans[8233]<=tmp[8132]*kernel[0]+tmp[8133]*kernel[1]+tmp[8134]*kernel[2]+tmp[8232]*kernel[3]+tmp[8233]*kernel[4]+tmp[8234]*kernel[5]+tmp[8332]*kernel[6]+tmp[8333]*kernel[7]+tmp[8334]*kernel[8];
				ans[8234]<=tmp[8133]*kernel[0]+tmp[8134]*kernel[1]+tmp[8135]*kernel[2]+tmp[8233]*kernel[3]+tmp[8234]*kernel[4]+tmp[8235]*kernel[5]+tmp[8333]*kernel[6]+tmp[8334]*kernel[7]+tmp[8335]*kernel[8];
				ans[8235]<=tmp[8134]*kernel[0]+tmp[8135]*kernel[1]+tmp[8136]*kernel[2]+tmp[8234]*kernel[3]+tmp[8235]*kernel[4]+tmp[8236]*kernel[5]+tmp[8334]*kernel[6]+tmp[8335]*kernel[7]+tmp[8336]*kernel[8];
				ans[8236]<=tmp[8135]*kernel[0]+tmp[8136]*kernel[1]+tmp[8137]*kernel[2]+tmp[8235]*kernel[3]+tmp[8236]*kernel[4]+tmp[8237]*kernel[5]+tmp[8335]*kernel[6]+tmp[8336]*kernel[7]+tmp[8337]*kernel[8];
				ans[8237]<=tmp[8136]*kernel[0]+tmp[8137]*kernel[1]+tmp[8138]*kernel[2]+tmp[8236]*kernel[3]+tmp[8237]*kernel[4]+tmp[8238]*kernel[5]+tmp[8336]*kernel[6]+tmp[8337]*kernel[7]+tmp[8338]*kernel[8];
				ans[8238]<=tmp[8137]*kernel[0]+tmp[8138]*kernel[1]+tmp[8139]*kernel[2]+tmp[8237]*kernel[3]+tmp[8238]*kernel[4]+tmp[8239]*kernel[5]+tmp[8337]*kernel[6]+tmp[8338]*kernel[7]+tmp[8339]*kernel[8];
				ans[8239]<=tmp[8138]*kernel[0]+tmp[8139]*kernel[1]+tmp[8140]*kernel[2]+tmp[8238]*kernel[3]+tmp[8239]*kernel[4]+tmp[8240]*kernel[5]+tmp[8338]*kernel[6]+tmp[8339]*kernel[7]+tmp[8340]*kernel[8];
				ans[8240]<=tmp[8139]*kernel[0]+tmp[8140]*kernel[1]+tmp[8141]*kernel[2]+tmp[8239]*kernel[3]+tmp[8240]*kernel[4]+tmp[8241]*kernel[5]+tmp[8339]*kernel[6]+tmp[8340]*kernel[7]+tmp[8341]*kernel[8];
				ans[8241]<=tmp[8140]*kernel[0]+tmp[8141]*kernel[1]+tmp[8142]*kernel[2]+tmp[8240]*kernel[3]+tmp[8241]*kernel[4]+tmp[8242]*kernel[5]+tmp[8340]*kernel[6]+tmp[8341]*kernel[7]+tmp[8342]*kernel[8];
				ans[8242]<=tmp[8141]*kernel[0]+tmp[8142]*kernel[1]+tmp[8143]*kernel[2]+tmp[8241]*kernel[3]+tmp[8242]*kernel[4]+tmp[8243]*kernel[5]+tmp[8341]*kernel[6]+tmp[8342]*kernel[7]+tmp[8343]*kernel[8];
				ans[8243]<=tmp[8142]*kernel[0]+tmp[8143]*kernel[1]+tmp[8144]*kernel[2]+tmp[8242]*kernel[3]+tmp[8243]*kernel[4]+tmp[8244]*kernel[5]+tmp[8342]*kernel[6]+tmp[8343]*kernel[7]+tmp[8344]*kernel[8];
				ans[8244]<=tmp[8143]*kernel[0]+tmp[8144]*kernel[1]+tmp[8145]*kernel[2]+tmp[8243]*kernel[3]+tmp[8244]*kernel[4]+tmp[8245]*kernel[5]+tmp[8343]*kernel[6]+tmp[8344]*kernel[7]+tmp[8345]*kernel[8];
				ans[8245]<=tmp[8144]*kernel[0]+tmp[8145]*kernel[1]+tmp[8146]*kernel[2]+tmp[8244]*kernel[3]+tmp[8245]*kernel[4]+tmp[8246]*kernel[5]+tmp[8344]*kernel[6]+tmp[8345]*kernel[7]+tmp[8346]*kernel[8];
				ans[8246]<=tmp[8145]*kernel[0]+tmp[8146]*kernel[1]+tmp[8147]*kernel[2]+tmp[8245]*kernel[3]+tmp[8246]*kernel[4]+tmp[8247]*kernel[5]+tmp[8345]*kernel[6]+tmp[8346]*kernel[7]+tmp[8347]*kernel[8];
				ans[8247]<=tmp[8146]*kernel[0]+tmp[8147]*kernel[1]+tmp[8148]*kernel[2]+tmp[8246]*kernel[3]+tmp[8247]*kernel[4]+tmp[8248]*kernel[5]+tmp[8346]*kernel[6]+tmp[8347]*kernel[7]+tmp[8348]*kernel[8];
				ans[8248]<=tmp[8147]*kernel[0]+tmp[8148]*kernel[1]+tmp[8149]*kernel[2]+tmp[8247]*kernel[3]+tmp[8248]*kernel[4]+tmp[8249]*kernel[5]+tmp[8347]*kernel[6]+tmp[8348]*kernel[7]+tmp[8349]*kernel[8];
				ans[8249]<=tmp[8148]*kernel[0]+tmp[8149]*kernel[1]+tmp[8150]*kernel[2]+tmp[8248]*kernel[3]+tmp[8249]*kernel[4]+tmp[8250]*kernel[5]+tmp[8348]*kernel[6]+tmp[8349]*kernel[7]+tmp[8350]*kernel[8];
				ans[8250]<=tmp[8149]*kernel[0]+tmp[8150]*kernel[1]+tmp[8151]*kernel[2]+tmp[8249]*kernel[3]+tmp[8250]*kernel[4]+tmp[8251]*kernel[5]+tmp[8349]*kernel[6]+tmp[8350]*kernel[7]+tmp[8351]*kernel[8];
				ans[8251]<=tmp[8150]*kernel[0]+tmp[8151]*kernel[1]+tmp[8152]*kernel[2]+tmp[8250]*kernel[3]+tmp[8251]*kernel[4]+tmp[8252]*kernel[5]+tmp[8350]*kernel[6]+tmp[8351]*kernel[7]+tmp[8352]*kernel[8];
				ans[8252]<=tmp[8151]*kernel[0]+tmp[8152]*kernel[1]+tmp[8153]*kernel[2]+tmp[8251]*kernel[3]+tmp[8252]*kernel[4]+tmp[8253]*kernel[5]+tmp[8351]*kernel[6]+tmp[8352]*kernel[7]+tmp[8353]*kernel[8];
				ans[8253]<=tmp[8152]*kernel[0]+tmp[8153]*kernel[1]+tmp[8154]*kernel[2]+tmp[8252]*kernel[3]+tmp[8253]*kernel[4]+tmp[8254]*kernel[5]+tmp[8352]*kernel[6]+tmp[8353]*kernel[7]+tmp[8354]*kernel[8];
				ans[8254]<=tmp[8153]*kernel[0]+tmp[8154]*kernel[1]+tmp[8155]*kernel[2]+tmp[8253]*kernel[3]+tmp[8254]*kernel[4]+tmp[8255]*kernel[5]+tmp[8353]*kernel[6]+tmp[8354]*kernel[7]+tmp[8355]*kernel[8];
				ans[8255]<=tmp[8154]*kernel[0]+tmp[8155]*kernel[1]+tmp[8156]*kernel[2]+tmp[8254]*kernel[3]+tmp[8255]*kernel[4]+tmp[8256]*kernel[5]+tmp[8354]*kernel[6]+tmp[8355]*kernel[7]+tmp[8356]*kernel[8];
				ans[8256]<=tmp[8155]*kernel[0]+tmp[8156]*kernel[1]+tmp[8157]*kernel[2]+tmp[8255]*kernel[3]+tmp[8256]*kernel[4]+tmp[8257]*kernel[5]+tmp[8355]*kernel[6]+tmp[8356]*kernel[7]+tmp[8357]*kernel[8];
				ans[8257]<=tmp[8156]*kernel[0]+tmp[8157]*kernel[1]+tmp[8158]*kernel[2]+tmp[8256]*kernel[3]+tmp[8257]*kernel[4]+tmp[8258]*kernel[5]+tmp[8356]*kernel[6]+tmp[8357]*kernel[7]+tmp[8358]*kernel[8];
				ans[8258]<=tmp[8157]*kernel[0]+tmp[8158]*kernel[1]+tmp[8159]*kernel[2]+tmp[8257]*kernel[3]+tmp[8258]*kernel[4]+tmp[8259]*kernel[5]+tmp[8357]*kernel[6]+tmp[8358]*kernel[7]+tmp[8359]*kernel[8];
				ans[8259]<=tmp[8158]*kernel[0]+tmp[8159]*kernel[1]+tmp[8160]*kernel[2]+tmp[8258]*kernel[3]+tmp[8259]*kernel[4]+tmp[8260]*kernel[5]+tmp[8358]*kernel[6]+tmp[8359]*kernel[7]+tmp[8360]*kernel[8];
				ans[8260]<=tmp[8159]*kernel[0]+tmp[8160]*kernel[1]+tmp[8161]*kernel[2]+tmp[8259]*kernel[3]+tmp[8260]*kernel[4]+tmp[8261]*kernel[5]+tmp[8359]*kernel[6]+tmp[8360]*kernel[7]+tmp[8361]*kernel[8];
				ans[8261]<=tmp[8160]*kernel[0]+tmp[8161]*kernel[1]+tmp[8162]*kernel[2]+tmp[8260]*kernel[3]+tmp[8261]*kernel[4]+tmp[8262]*kernel[5]+tmp[8360]*kernel[6]+tmp[8361]*kernel[7]+tmp[8362]*kernel[8];
				ans[8262]<=tmp[8161]*kernel[0]+tmp[8162]*kernel[1]+tmp[8163]*kernel[2]+tmp[8261]*kernel[3]+tmp[8262]*kernel[4]+tmp[8263]*kernel[5]+tmp[8361]*kernel[6]+tmp[8362]*kernel[7]+tmp[8363]*kernel[8];
				ans[8263]<=tmp[8162]*kernel[0]+tmp[8163]*kernel[1]+tmp[8164]*kernel[2]+tmp[8262]*kernel[3]+tmp[8263]*kernel[4]+tmp[8264]*kernel[5]+tmp[8362]*kernel[6]+tmp[8363]*kernel[7]+tmp[8364]*kernel[8];
				ans[8264]<=tmp[8163]*kernel[0]+tmp[8164]*kernel[1]+tmp[8165]*kernel[2]+tmp[8263]*kernel[3]+tmp[8264]*kernel[4]+tmp[8265]*kernel[5]+tmp[8363]*kernel[6]+tmp[8364]*kernel[7]+tmp[8365]*kernel[8];
				ans[8265]<=tmp[8164]*kernel[0]+tmp[8165]*kernel[1]+tmp[8166]*kernel[2]+tmp[8264]*kernel[3]+tmp[8265]*kernel[4]+tmp[8266]*kernel[5]+tmp[8364]*kernel[6]+tmp[8365]*kernel[7]+tmp[8366]*kernel[8];
				ans[8266]<=tmp[8165]*kernel[0]+tmp[8166]*kernel[1]+tmp[8167]*kernel[2]+tmp[8265]*kernel[3]+tmp[8266]*kernel[4]+tmp[8267]*kernel[5]+tmp[8365]*kernel[6]+tmp[8366]*kernel[7]+tmp[8367]*kernel[8];
				ans[8267]<=tmp[8166]*kernel[0]+tmp[8167]*kernel[1]+tmp[8168]*kernel[2]+tmp[8266]*kernel[3]+tmp[8267]*kernel[4]+tmp[8268]*kernel[5]+tmp[8366]*kernel[6]+tmp[8367]*kernel[7]+tmp[8368]*kernel[8];
				ans[8268]<=tmp[8167]*kernel[0]+tmp[8168]*kernel[1]+tmp[8169]*kernel[2]+tmp[8267]*kernel[3]+tmp[8268]*kernel[4]+tmp[8269]*kernel[5]+tmp[8367]*kernel[6]+tmp[8368]*kernel[7]+tmp[8369]*kernel[8];
				ans[8269]<=tmp[8168]*kernel[0]+tmp[8169]*kernel[1]+tmp[8170]*kernel[2]+tmp[8268]*kernel[3]+tmp[8269]*kernel[4]+tmp[8270]*kernel[5]+tmp[8368]*kernel[6]+tmp[8369]*kernel[7]+tmp[8370]*kernel[8];
				ans[8270]<=tmp[8169]*kernel[0]+tmp[8170]*kernel[1]+tmp[8171]*kernel[2]+tmp[8269]*kernel[3]+tmp[8270]*kernel[4]+tmp[8271]*kernel[5]+tmp[8369]*kernel[6]+tmp[8370]*kernel[7]+tmp[8371]*kernel[8];
				ans[8271]<=tmp[8170]*kernel[0]+tmp[8171]*kernel[1]+tmp[8172]*kernel[2]+tmp[8270]*kernel[3]+tmp[8271]*kernel[4]+tmp[8272]*kernel[5]+tmp[8370]*kernel[6]+tmp[8371]*kernel[7]+tmp[8372]*kernel[8];
				ans[8272]<=tmp[8171]*kernel[0]+tmp[8172]*kernel[1]+tmp[8173]*kernel[2]+tmp[8271]*kernel[3]+tmp[8272]*kernel[4]+tmp[8273]*kernel[5]+tmp[8371]*kernel[6]+tmp[8372]*kernel[7]+tmp[8373]*kernel[8];
				ans[8273]<=tmp[8172]*kernel[0]+tmp[8173]*kernel[1]+tmp[8174]*kernel[2]+tmp[8272]*kernel[3]+tmp[8273]*kernel[4]+tmp[8274]*kernel[5]+tmp[8372]*kernel[6]+tmp[8373]*kernel[7]+tmp[8374]*kernel[8];
				ans[8274]<=tmp[8173]*kernel[0]+tmp[8174]*kernel[1]+tmp[8175]*kernel[2]+tmp[8273]*kernel[3]+tmp[8274]*kernel[4]+tmp[8275]*kernel[5]+tmp[8373]*kernel[6]+tmp[8374]*kernel[7]+tmp[8375]*kernel[8];
				ans[8275]<=tmp[8174]*kernel[0]+tmp[8175]*kernel[1]+tmp[8176]*kernel[2]+tmp[8274]*kernel[3]+tmp[8275]*kernel[4]+tmp[8276]*kernel[5]+tmp[8374]*kernel[6]+tmp[8375]*kernel[7]+tmp[8376]*kernel[8];
				ans[8276]<=tmp[8175]*kernel[0]+tmp[8176]*kernel[1]+tmp[8177]*kernel[2]+tmp[8275]*kernel[3]+tmp[8276]*kernel[4]+tmp[8277]*kernel[5]+tmp[8375]*kernel[6]+tmp[8376]*kernel[7]+tmp[8377]*kernel[8];
				ans[8277]<=tmp[8176]*kernel[0]+tmp[8177]*kernel[1]+tmp[8178]*kernel[2]+tmp[8276]*kernel[3]+tmp[8277]*kernel[4]+tmp[8278]*kernel[5]+tmp[8376]*kernel[6]+tmp[8377]*kernel[7]+tmp[8378]*kernel[8];
				ans[8278]<=tmp[8177]*kernel[0]+tmp[8178]*kernel[1]+tmp[8179]*kernel[2]+tmp[8277]*kernel[3]+tmp[8278]*kernel[4]+tmp[8279]*kernel[5]+tmp[8377]*kernel[6]+tmp[8378]*kernel[7]+tmp[8379]*kernel[8];
				ans[8279]<=tmp[8178]*kernel[0]+tmp[8179]*kernel[1]+tmp[8180]*kernel[2]+tmp[8278]*kernel[3]+tmp[8279]*kernel[4]+tmp[8280]*kernel[5]+tmp[8378]*kernel[6]+tmp[8379]*kernel[7]+tmp[8380]*kernel[8];
				ans[8280]<=tmp[8179]*kernel[0]+tmp[8180]*kernel[1]+tmp[8181]*kernel[2]+tmp[8279]*kernel[3]+tmp[8280]*kernel[4]+tmp[8281]*kernel[5]+tmp[8379]*kernel[6]+tmp[8380]*kernel[7]+tmp[8381]*kernel[8];
				ans[8281]<=tmp[8180]*kernel[0]+tmp[8181]*kernel[1]+tmp[8182]*kernel[2]+tmp[8280]*kernel[3]+tmp[8281]*kernel[4]+tmp[8282]*kernel[5]+tmp[8380]*kernel[6]+tmp[8381]*kernel[7]+tmp[8382]*kernel[8];
				ans[8282]<=tmp[8181]*kernel[0]+tmp[8182]*kernel[1]+tmp[8183]*kernel[2]+tmp[8281]*kernel[3]+tmp[8282]*kernel[4]+tmp[8283]*kernel[5]+tmp[8381]*kernel[6]+tmp[8382]*kernel[7]+tmp[8383]*kernel[8];
				ans[8283]<=tmp[8182]*kernel[0]+tmp[8183]*kernel[1]+tmp[8184]*kernel[2]+tmp[8282]*kernel[3]+tmp[8283]*kernel[4]+tmp[8284]*kernel[5]+tmp[8382]*kernel[6]+tmp[8383]*kernel[7]+tmp[8384]*kernel[8];
				ans[8284]<=tmp[8183]*kernel[0]+tmp[8184]*kernel[1]+tmp[8185]*kernel[2]+tmp[8283]*kernel[3]+tmp[8284]*kernel[4]+tmp[8285]*kernel[5]+tmp[8383]*kernel[6]+tmp[8384]*kernel[7]+tmp[8385]*kernel[8];
				ans[8285]<=tmp[8184]*kernel[0]+tmp[8185]*kernel[1]+tmp[8186]*kernel[2]+tmp[8284]*kernel[3]+tmp[8285]*kernel[4]+tmp[8286]*kernel[5]+tmp[8384]*kernel[6]+tmp[8385]*kernel[7]+tmp[8386]*kernel[8];
				ans[8286]<=tmp[8185]*kernel[0]+tmp[8186]*kernel[1]+tmp[8187]*kernel[2]+tmp[8285]*kernel[3]+tmp[8286]*kernel[4]+tmp[8287]*kernel[5]+tmp[8385]*kernel[6]+tmp[8386]*kernel[7]+tmp[8387]*kernel[8];
				ans[8287]<=tmp[8186]*kernel[0]+tmp[8187]*kernel[1]+tmp[8188]*kernel[2]+tmp[8286]*kernel[3]+tmp[8287]*kernel[4]+tmp[8288]*kernel[5]+tmp[8386]*kernel[6]+tmp[8387]*kernel[7]+tmp[8388]*kernel[8];
				ans[8288]<=tmp[8187]*kernel[0]+tmp[8188]*kernel[1]+tmp[8189]*kernel[2]+tmp[8287]*kernel[3]+tmp[8288]*kernel[4]+tmp[8289]*kernel[5]+tmp[8387]*kernel[6]+tmp[8388]*kernel[7]+tmp[8389]*kernel[8];
				ans[8289]<=tmp[8188]*kernel[0]+tmp[8189]*kernel[1]+tmp[8190]*kernel[2]+tmp[8288]*kernel[3]+tmp[8289]*kernel[4]+tmp[8290]*kernel[5]+tmp[8388]*kernel[6]+tmp[8389]*kernel[7]+tmp[8390]*kernel[8];
				ans[8290]<=tmp[8189]*kernel[0]+tmp[8190]*kernel[1]+tmp[8191]*kernel[2]+tmp[8289]*kernel[3]+tmp[8290]*kernel[4]+tmp[8291]*kernel[5]+tmp[8389]*kernel[6]+tmp[8390]*kernel[7]+tmp[8391]*kernel[8];
				ans[8291]<=tmp[8190]*kernel[0]+tmp[8191]*kernel[1]+tmp[8192]*kernel[2]+tmp[8290]*kernel[3]+tmp[8291]*kernel[4]+tmp[8292]*kernel[5]+tmp[8390]*kernel[6]+tmp[8391]*kernel[7]+tmp[8392]*kernel[8];
				ans[8292]<=tmp[8191]*kernel[0]+tmp[8192]*kernel[1]+tmp[8193]*kernel[2]+tmp[8291]*kernel[3]+tmp[8292]*kernel[4]+tmp[8293]*kernel[5]+tmp[8391]*kernel[6]+tmp[8392]*kernel[7]+tmp[8393]*kernel[8];
				ans[8293]<=tmp[8192]*kernel[0]+tmp[8193]*kernel[1]+tmp[8194]*kernel[2]+tmp[8292]*kernel[3]+tmp[8293]*kernel[4]+tmp[8294]*kernel[5]+tmp[8392]*kernel[6]+tmp[8393]*kernel[7]+tmp[8394]*kernel[8];
				ans[8294]<=tmp[8193]*kernel[0]+tmp[8194]*kernel[1]+tmp[8195]*kernel[2]+tmp[8293]*kernel[3]+tmp[8294]*kernel[4]+tmp[8295]*kernel[5]+tmp[8393]*kernel[6]+tmp[8394]*kernel[7]+tmp[8395]*kernel[8];
				ans[8295]<=tmp[8194]*kernel[0]+tmp[8195]*kernel[1]+tmp[8196]*kernel[2]+tmp[8294]*kernel[3]+tmp[8295]*kernel[4]+tmp[8296]*kernel[5]+tmp[8394]*kernel[6]+tmp[8395]*kernel[7]+tmp[8396]*kernel[8];
				ans[8296]<=tmp[8195]*kernel[0]+tmp[8196]*kernel[1]+tmp[8197]*kernel[2]+tmp[8295]*kernel[3]+tmp[8296]*kernel[4]+tmp[8297]*kernel[5]+tmp[8395]*kernel[6]+tmp[8396]*kernel[7]+tmp[8397]*kernel[8];
				ans[8297]<=tmp[8196]*kernel[0]+tmp[8197]*kernel[1]+tmp[8198]*kernel[2]+tmp[8296]*kernel[3]+tmp[8297]*kernel[4]+tmp[8298]*kernel[5]+tmp[8396]*kernel[6]+tmp[8397]*kernel[7]+tmp[8398]*kernel[8];
				ans[8298]<=tmp[8197]*kernel[0]+tmp[8198]*kernel[1]+tmp[8199]*kernel[2]+tmp[8297]*kernel[3]+tmp[8298]*kernel[4]+tmp[8299]*kernel[5]+tmp[8397]*kernel[6]+tmp[8398]*kernel[7]+tmp[8399]*kernel[8];
				ans[8299]<=tmp[8198]*kernel[0]+tmp[8199]*kernel[1]+tmp[8298]*kernel[3]+tmp[8299]*kernel[4]+tmp[8398]*kernel[6]+tmp[8399]*kernel[7];
				ans[8300]<=tmp[8200]*kernel[1]+tmp[8201]*kernel[2]+tmp[8300]*kernel[4]+tmp[8301]*kernel[5]+tmp[8400]*kernel[7]+tmp[8401]*kernel[8];
				ans[8301]<=tmp[8200]*kernel[0]+tmp[8201]*kernel[1]+tmp[8202]*kernel[2]+tmp[8300]*kernel[3]+tmp[8301]*kernel[4]+tmp[8302]*kernel[5]+tmp[8400]*kernel[6]+tmp[8401]*kernel[7]+tmp[8402]*kernel[8];
				ans[8302]<=tmp[8201]*kernel[0]+tmp[8202]*kernel[1]+tmp[8203]*kernel[2]+tmp[8301]*kernel[3]+tmp[8302]*kernel[4]+tmp[8303]*kernel[5]+tmp[8401]*kernel[6]+tmp[8402]*kernel[7]+tmp[8403]*kernel[8];
				ans[8303]<=tmp[8202]*kernel[0]+tmp[8203]*kernel[1]+tmp[8204]*kernel[2]+tmp[8302]*kernel[3]+tmp[8303]*kernel[4]+tmp[8304]*kernel[5]+tmp[8402]*kernel[6]+tmp[8403]*kernel[7]+tmp[8404]*kernel[8];
				ans[8304]<=tmp[8203]*kernel[0]+tmp[8204]*kernel[1]+tmp[8205]*kernel[2]+tmp[8303]*kernel[3]+tmp[8304]*kernel[4]+tmp[8305]*kernel[5]+tmp[8403]*kernel[6]+tmp[8404]*kernel[7]+tmp[8405]*kernel[8];
				ans[8305]<=tmp[8204]*kernel[0]+tmp[8205]*kernel[1]+tmp[8206]*kernel[2]+tmp[8304]*kernel[3]+tmp[8305]*kernel[4]+tmp[8306]*kernel[5]+tmp[8404]*kernel[6]+tmp[8405]*kernel[7]+tmp[8406]*kernel[8];
				ans[8306]<=tmp[8205]*kernel[0]+tmp[8206]*kernel[1]+tmp[8207]*kernel[2]+tmp[8305]*kernel[3]+tmp[8306]*kernel[4]+tmp[8307]*kernel[5]+tmp[8405]*kernel[6]+tmp[8406]*kernel[7]+tmp[8407]*kernel[8];
				ans[8307]<=tmp[8206]*kernel[0]+tmp[8207]*kernel[1]+tmp[8208]*kernel[2]+tmp[8306]*kernel[3]+tmp[8307]*kernel[4]+tmp[8308]*kernel[5]+tmp[8406]*kernel[6]+tmp[8407]*kernel[7]+tmp[8408]*kernel[8];
				ans[8308]<=tmp[8207]*kernel[0]+tmp[8208]*kernel[1]+tmp[8209]*kernel[2]+tmp[8307]*kernel[3]+tmp[8308]*kernel[4]+tmp[8309]*kernel[5]+tmp[8407]*kernel[6]+tmp[8408]*kernel[7]+tmp[8409]*kernel[8];
				ans[8309]<=tmp[8208]*kernel[0]+tmp[8209]*kernel[1]+tmp[8210]*kernel[2]+tmp[8308]*kernel[3]+tmp[8309]*kernel[4]+tmp[8310]*kernel[5]+tmp[8408]*kernel[6]+tmp[8409]*kernel[7]+tmp[8410]*kernel[8];
				ans[8310]<=tmp[8209]*kernel[0]+tmp[8210]*kernel[1]+tmp[8211]*kernel[2]+tmp[8309]*kernel[3]+tmp[8310]*kernel[4]+tmp[8311]*kernel[5]+tmp[8409]*kernel[6]+tmp[8410]*kernel[7]+tmp[8411]*kernel[8];
				ans[8311]<=tmp[8210]*kernel[0]+tmp[8211]*kernel[1]+tmp[8212]*kernel[2]+tmp[8310]*kernel[3]+tmp[8311]*kernel[4]+tmp[8312]*kernel[5]+tmp[8410]*kernel[6]+tmp[8411]*kernel[7]+tmp[8412]*kernel[8];
				ans[8312]<=tmp[8211]*kernel[0]+tmp[8212]*kernel[1]+tmp[8213]*kernel[2]+tmp[8311]*kernel[3]+tmp[8312]*kernel[4]+tmp[8313]*kernel[5]+tmp[8411]*kernel[6]+tmp[8412]*kernel[7]+tmp[8413]*kernel[8];
				ans[8313]<=tmp[8212]*kernel[0]+tmp[8213]*kernel[1]+tmp[8214]*kernel[2]+tmp[8312]*kernel[3]+tmp[8313]*kernel[4]+tmp[8314]*kernel[5]+tmp[8412]*kernel[6]+tmp[8413]*kernel[7]+tmp[8414]*kernel[8];
				ans[8314]<=tmp[8213]*kernel[0]+tmp[8214]*kernel[1]+tmp[8215]*kernel[2]+tmp[8313]*kernel[3]+tmp[8314]*kernel[4]+tmp[8315]*kernel[5]+tmp[8413]*kernel[6]+tmp[8414]*kernel[7]+tmp[8415]*kernel[8];
				ans[8315]<=tmp[8214]*kernel[0]+tmp[8215]*kernel[1]+tmp[8216]*kernel[2]+tmp[8314]*kernel[3]+tmp[8315]*kernel[4]+tmp[8316]*kernel[5]+tmp[8414]*kernel[6]+tmp[8415]*kernel[7]+tmp[8416]*kernel[8];
				ans[8316]<=tmp[8215]*kernel[0]+tmp[8216]*kernel[1]+tmp[8217]*kernel[2]+tmp[8315]*kernel[3]+tmp[8316]*kernel[4]+tmp[8317]*kernel[5]+tmp[8415]*kernel[6]+tmp[8416]*kernel[7]+tmp[8417]*kernel[8];
				ans[8317]<=tmp[8216]*kernel[0]+tmp[8217]*kernel[1]+tmp[8218]*kernel[2]+tmp[8316]*kernel[3]+tmp[8317]*kernel[4]+tmp[8318]*kernel[5]+tmp[8416]*kernel[6]+tmp[8417]*kernel[7]+tmp[8418]*kernel[8];
				ans[8318]<=tmp[8217]*kernel[0]+tmp[8218]*kernel[1]+tmp[8219]*kernel[2]+tmp[8317]*kernel[3]+tmp[8318]*kernel[4]+tmp[8319]*kernel[5]+tmp[8417]*kernel[6]+tmp[8418]*kernel[7]+tmp[8419]*kernel[8];
				ans[8319]<=tmp[8218]*kernel[0]+tmp[8219]*kernel[1]+tmp[8220]*kernel[2]+tmp[8318]*kernel[3]+tmp[8319]*kernel[4]+tmp[8320]*kernel[5]+tmp[8418]*kernel[6]+tmp[8419]*kernel[7]+tmp[8420]*kernel[8];
				ans[8320]<=tmp[8219]*kernel[0]+tmp[8220]*kernel[1]+tmp[8221]*kernel[2]+tmp[8319]*kernel[3]+tmp[8320]*kernel[4]+tmp[8321]*kernel[5]+tmp[8419]*kernel[6]+tmp[8420]*kernel[7]+tmp[8421]*kernel[8];
				ans[8321]<=tmp[8220]*kernel[0]+tmp[8221]*kernel[1]+tmp[8222]*kernel[2]+tmp[8320]*kernel[3]+tmp[8321]*kernel[4]+tmp[8322]*kernel[5]+tmp[8420]*kernel[6]+tmp[8421]*kernel[7]+tmp[8422]*kernel[8];
				ans[8322]<=tmp[8221]*kernel[0]+tmp[8222]*kernel[1]+tmp[8223]*kernel[2]+tmp[8321]*kernel[3]+tmp[8322]*kernel[4]+tmp[8323]*kernel[5]+tmp[8421]*kernel[6]+tmp[8422]*kernel[7]+tmp[8423]*kernel[8];
				ans[8323]<=tmp[8222]*kernel[0]+tmp[8223]*kernel[1]+tmp[8224]*kernel[2]+tmp[8322]*kernel[3]+tmp[8323]*kernel[4]+tmp[8324]*kernel[5]+tmp[8422]*kernel[6]+tmp[8423]*kernel[7]+tmp[8424]*kernel[8];
				ans[8324]<=tmp[8223]*kernel[0]+tmp[8224]*kernel[1]+tmp[8225]*kernel[2]+tmp[8323]*kernel[3]+tmp[8324]*kernel[4]+tmp[8325]*kernel[5]+tmp[8423]*kernel[6]+tmp[8424]*kernel[7]+tmp[8425]*kernel[8];
				ans[8325]<=tmp[8224]*kernel[0]+tmp[8225]*kernel[1]+tmp[8226]*kernel[2]+tmp[8324]*kernel[3]+tmp[8325]*kernel[4]+tmp[8326]*kernel[5]+tmp[8424]*kernel[6]+tmp[8425]*kernel[7]+tmp[8426]*kernel[8];
				ans[8326]<=tmp[8225]*kernel[0]+tmp[8226]*kernel[1]+tmp[8227]*kernel[2]+tmp[8325]*kernel[3]+tmp[8326]*kernel[4]+tmp[8327]*kernel[5]+tmp[8425]*kernel[6]+tmp[8426]*kernel[7]+tmp[8427]*kernel[8];
				ans[8327]<=tmp[8226]*kernel[0]+tmp[8227]*kernel[1]+tmp[8228]*kernel[2]+tmp[8326]*kernel[3]+tmp[8327]*kernel[4]+tmp[8328]*kernel[5]+tmp[8426]*kernel[6]+tmp[8427]*kernel[7]+tmp[8428]*kernel[8];
				ans[8328]<=tmp[8227]*kernel[0]+tmp[8228]*kernel[1]+tmp[8229]*kernel[2]+tmp[8327]*kernel[3]+tmp[8328]*kernel[4]+tmp[8329]*kernel[5]+tmp[8427]*kernel[6]+tmp[8428]*kernel[7]+tmp[8429]*kernel[8];
				ans[8329]<=tmp[8228]*kernel[0]+tmp[8229]*kernel[1]+tmp[8230]*kernel[2]+tmp[8328]*kernel[3]+tmp[8329]*kernel[4]+tmp[8330]*kernel[5]+tmp[8428]*kernel[6]+tmp[8429]*kernel[7]+tmp[8430]*kernel[8];
				ans[8330]<=tmp[8229]*kernel[0]+tmp[8230]*kernel[1]+tmp[8231]*kernel[2]+tmp[8329]*kernel[3]+tmp[8330]*kernel[4]+tmp[8331]*kernel[5]+tmp[8429]*kernel[6]+tmp[8430]*kernel[7]+tmp[8431]*kernel[8];
				ans[8331]<=tmp[8230]*kernel[0]+tmp[8231]*kernel[1]+tmp[8232]*kernel[2]+tmp[8330]*kernel[3]+tmp[8331]*kernel[4]+tmp[8332]*kernel[5]+tmp[8430]*kernel[6]+tmp[8431]*kernel[7]+tmp[8432]*kernel[8];
				ans[8332]<=tmp[8231]*kernel[0]+tmp[8232]*kernel[1]+tmp[8233]*kernel[2]+tmp[8331]*kernel[3]+tmp[8332]*kernel[4]+tmp[8333]*kernel[5]+tmp[8431]*kernel[6]+tmp[8432]*kernel[7]+tmp[8433]*kernel[8];
				ans[8333]<=tmp[8232]*kernel[0]+tmp[8233]*kernel[1]+tmp[8234]*kernel[2]+tmp[8332]*kernel[3]+tmp[8333]*kernel[4]+tmp[8334]*kernel[5]+tmp[8432]*kernel[6]+tmp[8433]*kernel[7]+tmp[8434]*kernel[8];
				ans[8334]<=tmp[8233]*kernel[0]+tmp[8234]*kernel[1]+tmp[8235]*kernel[2]+tmp[8333]*kernel[3]+tmp[8334]*kernel[4]+tmp[8335]*kernel[5]+tmp[8433]*kernel[6]+tmp[8434]*kernel[7]+tmp[8435]*kernel[8];
				ans[8335]<=tmp[8234]*kernel[0]+tmp[8235]*kernel[1]+tmp[8236]*kernel[2]+tmp[8334]*kernel[3]+tmp[8335]*kernel[4]+tmp[8336]*kernel[5]+tmp[8434]*kernel[6]+tmp[8435]*kernel[7]+tmp[8436]*kernel[8];
				ans[8336]<=tmp[8235]*kernel[0]+tmp[8236]*kernel[1]+tmp[8237]*kernel[2]+tmp[8335]*kernel[3]+tmp[8336]*kernel[4]+tmp[8337]*kernel[5]+tmp[8435]*kernel[6]+tmp[8436]*kernel[7]+tmp[8437]*kernel[8];
				ans[8337]<=tmp[8236]*kernel[0]+tmp[8237]*kernel[1]+tmp[8238]*kernel[2]+tmp[8336]*kernel[3]+tmp[8337]*kernel[4]+tmp[8338]*kernel[5]+tmp[8436]*kernel[6]+tmp[8437]*kernel[7]+tmp[8438]*kernel[8];
				ans[8338]<=tmp[8237]*kernel[0]+tmp[8238]*kernel[1]+tmp[8239]*kernel[2]+tmp[8337]*kernel[3]+tmp[8338]*kernel[4]+tmp[8339]*kernel[5]+tmp[8437]*kernel[6]+tmp[8438]*kernel[7]+tmp[8439]*kernel[8];
				ans[8339]<=tmp[8238]*kernel[0]+tmp[8239]*kernel[1]+tmp[8240]*kernel[2]+tmp[8338]*kernel[3]+tmp[8339]*kernel[4]+tmp[8340]*kernel[5]+tmp[8438]*kernel[6]+tmp[8439]*kernel[7]+tmp[8440]*kernel[8];
				ans[8340]<=tmp[8239]*kernel[0]+tmp[8240]*kernel[1]+tmp[8241]*kernel[2]+tmp[8339]*kernel[3]+tmp[8340]*kernel[4]+tmp[8341]*kernel[5]+tmp[8439]*kernel[6]+tmp[8440]*kernel[7]+tmp[8441]*kernel[8];
				ans[8341]<=tmp[8240]*kernel[0]+tmp[8241]*kernel[1]+tmp[8242]*kernel[2]+tmp[8340]*kernel[3]+tmp[8341]*kernel[4]+tmp[8342]*kernel[5]+tmp[8440]*kernel[6]+tmp[8441]*kernel[7]+tmp[8442]*kernel[8];
				ans[8342]<=tmp[8241]*kernel[0]+tmp[8242]*kernel[1]+tmp[8243]*kernel[2]+tmp[8341]*kernel[3]+tmp[8342]*kernel[4]+tmp[8343]*kernel[5]+tmp[8441]*kernel[6]+tmp[8442]*kernel[7]+tmp[8443]*kernel[8];
				ans[8343]<=tmp[8242]*kernel[0]+tmp[8243]*kernel[1]+tmp[8244]*kernel[2]+tmp[8342]*kernel[3]+tmp[8343]*kernel[4]+tmp[8344]*kernel[5]+tmp[8442]*kernel[6]+tmp[8443]*kernel[7]+tmp[8444]*kernel[8];
				ans[8344]<=tmp[8243]*kernel[0]+tmp[8244]*kernel[1]+tmp[8245]*kernel[2]+tmp[8343]*kernel[3]+tmp[8344]*kernel[4]+tmp[8345]*kernel[5]+tmp[8443]*kernel[6]+tmp[8444]*kernel[7]+tmp[8445]*kernel[8];
				ans[8345]<=tmp[8244]*kernel[0]+tmp[8245]*kernel[1]+tmp[8246]*kernel[2]+tmp[8344]*kernel[3]+tmp[8345]*kernel[4]+tmp[8346]*kernel[5]+tmp[8444]*kernel[6]+tmp[8445]*kernel[7]+tmp[8446]*kernel[8];
				ans[8346]<=tmp[8245]*kernel[0]+tmp[8246]*kernel[1]+tmp[8247]*kernel[2]+tmp[8345]*kernel[3]+tmp[8346]*kernel[4]+tmp[8347]*kernel[5]+tmp[8445]*kernel[6]+tmp[8446]*kernel[7]+tmp[8447]*kernel[8];
				ans[8347]<=tmp[8246]*kernel[0]+tmp[8247]*kernel[1]+tmp[8248]*kernel[2]+tmp[8346]*kernel[3]+tmp[8347]*kernel[4]+tmp[8348]*kernel[5]+tmp[8446]*kernel[6]+tmp[8447]*kernel[7]+tmp[8448]*kernel[8];
				ans[8348]<=tmp[8247]*kernel[0]+tmp[8248]*kernel[1]+tmp[8249]*kernel[2]+tmp[8347]*kernel[3]+tmp[8348]*kernel[4]+tmp[8349]*kernel[5]+tmp[8447]*kernel[6]+tmp[8448]*kernel[7]+tmp[8449]*kernel[8];
				ans[8349]<=tmp[8248]*kernel[0]+tmp[8249]*kernel[1]+tmp[8250]*kernel[2]+tmp[8348]*kernel[3]+tmp[8349]*kernel[4]+tmp[8350]*kernel[5]+tmp[8448]*kernel[6]+tmp[8449]*kernel[7]+tmp[8450]*kernel[8];
				ans[8350]<=tmp[8249]*kernel[0]+tmp[8250]*kernel[1]+tmp[8251]*kernel[2]+tmp[8349]*kernel[3]+tmp[8350]*kernel[4]+tmp[8351]*kernel[5]+tmp[8449]*kernel[6]+tmp[8450]*kernel[7]+tmp[8451]*kernel[8];
				ans[8351]<=tmp[8250]*kernel[0]+tmp[8251]*kernel[1]+tmp[8252]*kernel[2]+tmp[8350]*kernel[3]+tmp[8351]*kernel[4]+tmp[8352]*kernel[5]+tmp[8450]*kernel[6]+tmp[8451]*kernel[7]+tmp[8452]*kernel[8];
				ans[8352]<=tmp[8251]*kernel[0]+tmp[8252]*kernel[1]+tmp[8253]*kernel[2]+tmp[8351]*kernel[3]+tmp[8352]*kernel[4]+tmp[8353]*kernel[5]+tmp[8451]*kernel[6]+tmp[8452]*kernel[7]+tmp[8453]*kernel[8];
				ans[8353]<=tmp[8252]*kernel[0]+tmp[8253]*kernel[1]+tmp[8254]*kernel[2]+tmp[8352]*kernel[3]+tmp[8353]*kernel[4]+tmp[8354]*kernel[5]+tmp[8452]*kernel[6]+tmp[8453]*kernel[7]+tmp[8454]*kernel[8];
				ans[8354]<=tmp[8253]*kernel[0]+tmp[8254]*kernel[1]+tmp[8255]*kernel[2]+tmp[8353]*kernel[3]+tmp[8354]*kernel[4]+tmp[8355]*kernel[5]+tmp[8453]*kernel[6]+tmp[8454]*kernel[7]+tmp[8455]*kernel[8];
				ans[8355]<=tmp[8254]*kernel[0]+tmp[8255]*kernel[1]+tmp[8256]*kernel[2]+tmp[8354]*kernel[3]+tmp[8355]*kernel[4]+tmp[8356]*kernel[5]+tmp[8454]*kernel[6]+tmp[8455]*kernel[7]+tmp[8456]*kernel[8];
				ans[8356]<=tmp[8255]*kernel[0]+tmp[8256]*kernel[1]+tmp[8257]*kernel[2]+tmp[8355]*kernel[3]+tmp[8356]*kernel[4]+tmp[8357]*kernel[5]+tmp[8455]*kernel[6]+tmp[8456]*kernel[7]+tmp[8457]*kernel[8];
				ans[8357]<=tmp[8256]*kernel[0]+tmp[8257]*kernel[1]+tmp[8258]*kernel[2]+tmp[8356]*kernel[3]+tmp[8357]*kernel[4]+tmp[8358]*kernel[5]+tmp[8456]*kernel[6]+tmp[8457]*kernel[7]+tmp[8458]*kernel[8];
				ans[8358]<=tmp[8257]*kernel[0]+tmp[8258]*kernel[1]+tmp[8259]*kernel[2]+tmp[8357]*kernel[3]+tmp[8358]*kernel[4]+tmp[8359]*kernel[5]+tmp[8457]*kernel[6]+tmp[8458]*kernel[7]+tmp[8459]*kernel[8];
				ans[8359]<=tmp[8258]*kernel[0]+tmp[8259]*kernel[1]+tmp[8260]*kernel[2]+tmp[8358]*kernel[3]+tmp[8359]*kernel[4]+tmp[8360]*kernel[5]+tmp[8458]*kernel[6]+tmp[8459]*kernel[7]+tmp[8460]*kernel[8];
				ans[8360]<=tmp[8259]*kernel[0]+tmp[8260]*kernel[1]+tmp[8261]*kernel[2]+tmp[8359]*kernel[3]+tmp[8360]*kernel[4]+tmp[8361]*kernel[5]+tmp[8459]*kernel[6]+tmp[8460]*kernel[7]+tmp[8461]*kernel[8];
				ans[8361]<=tmp[8260]*kernel[0]+tmp[8261]*kernel[1]+tmp[8262]*kernel[2]+tmp[8360]*kernel[3]+tmp[8361]*kernel[4]+tmp[8362]*kernel[5]+tmp[8460]*kernel[6]+tmp[8461]*kernel[7]+tmp[8462]*kernel[8];
				ans[8362]<=tmp[8261]*kernel[0]+tmp[8262]*kernel[1]+tmp[8263]*kernel[2]+tmp[8361]*kernel[3]+tmp[8362]*kernel[4]+tmp[8363]*kernel[5]+tmp[8461]*kernel[6]+tmp[8462]*kernel[7]+tmp[8463]*kernel[8];
				ans[8363]<=tmp[8262]*kernel[0]+tmp[8263]*kernel[1]+tmp[8264]*kernel[2]+tmp[8362]*kernel[3]+tmp[8363]*kernel[4]+tmp[8364]*kernel[5]+tmp[8462]*kernel[6]+tmp[8463]*kernel[7]+tmp[8464]*kernel[8];
				ans[8364]<=tmp[8263]*kernel[0]+tmp[8264]*kernel[1]+tmp[8265]*kernel[2]+tmp[8363]*kernel[3]+tmp[8364]*kernel[4]+tmp[8365]*kernel[5]+tmp[8463]*kernel[6]+tmp[8464]*kernel[7]+tmp[8465]*kernel[8];
				ans[8365]<=tmp[8264]*kernel[0]+tmp[8265]*kernel[1]+tmp[8266]*kernel[2]+tmp[8364]*kernel[3]+tmp[8365]*kernel[4]+tmp[8366]*kernel[5]+tmp[8464]*kernel[6]+tmp[8465]*kernel[7]+tmp[8466]*kernel[8];
				ans[8366]<=tmp[8265]*kernel[0]+tmp[8266]*kernel[1]+tmp[8267]*kernel[2]+tmp[8365]*kernel[3]+tmp[8366]*kernel[4]+tmp[8367]*kernel[5]+tmp[8465]*kernel[6]+tmp[8466]*kernel[7]+tmp[8467]*kernel[8];
				ans[8367]<=tmp[8266]*kernel[0]+tmp[8267]*kernel[1]+tmp[8268]*kernel[2]+tmp[8366]*kernel[3]+tmp[8367]*kernel[4]+tmp[8368]*kernel[5]+tmp[8466]*kernel[6]+tmp[8467]*kernel[7]+tmp[8468]*kernel[8];
				ans[8368]<=tmp[8267]*kernel[0]+tmp[8268]*kernel[1]+tmp[8269]*kernel[2]+tmp[8367]*kernel[3]+tmp[8368]*kernel[4]+tmp[8369]*kernel[5]+tmp[8467]*kernel[6]+tmp[8468]*kernel[7]+tmp[8469]*kernel[8];
				ans[8369]<=tmp[8268]*kernel[0]+tmp[8269]*kernel[1]+tmp[8270]*kernel[2]+tmp[8368]*kernel[3]+tmp[8369]*kernel[4]+tmp[8370]*kernel[5]+tmp[8468]*kernel[6]+tmp[8469]*kernel[7]+tmp[8470]*kernel[8];
				ans[8370]<=tmp[8269]*kernel[0]+tmp[8270]*kernel[1]+tmp[8271]*kernel[2]+tmp[8369]*kernel[3]+tmp[8370]*kernel[4]+tmp[8371]*kernel[5]+tmp[8469]*kernel[6]+tmp[8470]*kernel[7]+tmp[8471]*kernel[8];
				ans[8371]<=tmp[8270]*kernel[0]+tmp[8271]*kernel[1]+tmp[8272]*kernel[2]+tmp[8370]*kernel[3]+tmp[8371]*kernel[4]+tmp[8372]*kernel[5]+tmp[8470]*kernel[6]+tmp[8471]*kernel[7]+tmp[8472]*kernel[8];
				ans[8372]<=tmp[8271]*kernel[0]+tmp[8272]*kernel[1]+tmp[8273]*kernel[2]+tmp[8371]*kernel[3]+tmp[8372]*kernel[4]+tmp[8373]*kernel[5]+tmp[8471]*kernel[6]+tmp[8472]*kernel[7]+tmp[8473]*kernel[8];
				ans[8373]<=tmp[8272]*kernel[0]+tmp[8273]*kernel[1]+tmp[8274]*kernel[2]+tmp[8372]*kernel[3]+tmp[8373]*kernel[4]+tmp[8374]*kernel[5]+tmp[8472]*kernel[6]+tmp[8473]*kernel[7]+tmp[8474]*kernel[8];
				ans[8374]<=tmp[8273]*kernel[0]+tmp[8274]*kernel[1]+tmp[8275]*kernel[2]+tmp[8373]*kernel[3]+tmp[8374]*kernel[4]+tmp[8375]*kernel[5]+tmp[8473]*kernel[6]+tmp[8474]*kernel[7]+tmp[8475]*kernel[8];
				ans[8375]<=tmp[8274]*kernel[0]+tmp[8275]*kernel[1]+tmp[8276]*kernel[2]+tmp[8374]*kernel[3]+tmp[8375]*kernel[4]+tmp[8376]*kernel[5]+tmp[8474]*kernel[6]+tmp[8475]*kernel[7]+tmp[8476]*kernel[8];
				ans[8376]<=tmp[8275]*kernel[0]+tmp[8276]*kernel[1]+tmp[8277]*kernel[2]+tmp[8375]*kernel[3]+tmp[8376]*kernel[4]+tmp[8377]*kernel[5]+tmp[8475]*kernel[6]+tmp[8476]*kernel[7]+tmp[8477]*kernel[8];
				ans[8377]<=tmp[8276]*kernel[0]+tmp[8277]*kernel[1]+tmp[8278]*kernel[2]+tmp[8376]*kernel[3]+tmp[8377]*kernel[4]+tmp[8378]*kernel[5]+tmp[8476]*kernel[6]+tmp[8477]*kernel[7]+tmp[8478]*kernel[8];
				ans[8378]<=tmp[8277]*kernel[0]+tmp[8278]*kernel[1]+tmp[8279]*kernel[2]+tmp[8377]*kernel[3]+tmp[8378]*kernel[4]+tmp[8379]*kernel[5]+tmp[8477]*kernel[6]+tmp[8478]*kernel[7]+tmp[8479]*kernel[8];
				ans[8379]<=tmp[8278]*kernel[0]+tmp[8279]*kernel[1]+tmp[8280]*kernel[2]+tmp[8378]*kernel[3]+tmp[8379]*kernel[4]+tmp[8380]*kernel[5]+tmp[8478]*kernel[6]+tmp[8479]*kernel[7]+tmp[8480]*kernel[8];
				ans[8380]<=tmp[8279]*kernel[0]+tmp[8280]*kernel[1]+tmp[8281]*kernel[2]+tmp[8379]*kernel[3]+tmp[8380]*kernel[4]+tmp[8381]*kernel[5]+tmp[8479]*kernel[6]+tmp[8480]*kernel[7]+tmp[8481]*kernel[8];
				ans[8381]<=tmp[8280]*kernel[0]+tmp[8281]*kernel[1]+tmp[8282]*kernel[2]+tmp[8380]*kernel[3]+tmp[8381]*kernel[4]+tmp[8382]*kernel[5]+tmp[8480]*kernel[6]+tmp[8481]*kernel[7]+tmp[8482]*kernel[8];
				ans[8382]<=tmp[8281]*kernel[0]+tmp[8282]*kernel[1]+tmp[8283]*kernel[2]+tmp[8381]*kernel[3]+tmp[8382]*kernel[4]+tmp[8383]*kernel[5]+tmp[8481]*kernel[6]+tmp[8482]*kernel[7]+tmp[8483]*kernel[8];
				ans[8383]<=tmp[8282]*kernel[0]+tmp[8283]*kernel[1]+tmp[8284]*kernel[2]+tmp[8382]*kernel[3]+tmp[8383]*kernel[4]+tmp[8384]*kernel[5]+tmp[8482]*kernel[6]+tmp[8483]*kernel[7]+tmp[8484]*kernel[8];
				ans[8384]<=tmp[8283]*kernel[0]+tmp[8284]*kernel[1]+tmp[8285]*kernel[2]+tmp[8383]*kernel[3]+tmp[8384]*kernel[4]+tmp[8385]*kernel[5]+tmp[8483]*kernel[6]+tmp[8484]*kernel[7]+tmp[8485]*kernel[8];
				ans[8385]<=tmp[8284]*kernel[0]+tmp[8285]*kernel[1]+tmp[8286]*kernel[2]+tmp[8384]*kernel[3]+tmp[8385]*kernel[4]+tmp[8386]*kernel[5]+tmp[8484]*kernel[6]+tmp[8485]*kernel[7]+tmp[8486]*kernel[8];
				ans[8386]<=tmp[8285]*kernel[0]+tmp[8286]*kernel[1]+tmp[8287]*kernel[2]+tmp[8385]*kernel[3]+tmp[8386]*kernel[4]+tmp[8387]*kernel[5]+tmp[8485]*kernel[6]+tmp[8486]*kernel[7]+tmp[8487]*kernel[8];
				ans[8387]<=tmp[8286]*kernel[0]+tmp[8287]*kernel[1]+tmp[8288]*kernel[2]+tmp[8386]*kernel[3]+tmp[8387]*kernel[4]+tmp[8388]*kernel[5]+tmp[8486]*kernel[6]+tmp[8487]*kernel[7]+tmp[8488]*kernel[8];
				ans[8388]<=tmp[8287]*kernel[0]+tmp[8288]*kernel[1]+tmp[8289]*kernel[2]+tmp[8387]*kernel[3]+tmp[8388]*kernel[4]+tmp[8389]*kernel[5]+tmp[8487]*kernel[6]+tmp[8488]*kernel[7]+tmp[8489]*kernel[8];
				ans[8389]<=tmp[8288]*kernel[0]+tmp[8289]*kernel[1]+tmp[8290]*kernel[2]+tmp[8388]*kernel[3]+tmp[8389]*kernel[4]+tmp[8390]*kernel[5]+tmp[8488]*kernel[6]+tmp[8489]*kernel[7]+tmp[8490]*kernel[8];
				ans[8390]<=tmp[8289]*kernel[0]+tmp[8290]*kernel[1]+tmp[8291]*kernel[2]+tmp[8389]*kernel[3]+tmp[8390]*kernel[4]+tmp[8391]*kernel[5]+tmp[8489]*kernel[6]+tmp[8490]*kernel[7]+tmp[8491]*kernel[8];
				ans[8391]<=tmp[8290]*kernel[0]+tmp[8291]*kernel[1]+tmp[8292]*kernel[2]+tmp[8390]*kernel[3]+tmp[8391]*kernel[4]+tmp[8392]*kernel[5]+tmp[8490]*kernel[6]+tmp[8491]*kernel[7]+tmp[8492]*kernel[8];
				ans[8392]<=tmp[8291]*kernel[0]+tmp[8292]*kernel[1]+tmp[8293]*kernel[2]+tmp[8391]*kernel[3]+tmp[8392]*kernel[4]+tmp[8393]*kernel[5]+tmp[8491]*kernel[6]+tmp[8492]*kernel[7]+tmp[8493]*kernel[8];
				ans[8393]<=tmp[8292]*kernel[0]+tmp[8293]*kernel[1]+tmp[8294]*kernel[2]+tmp[8392]*kernel[3]+tmp[8393]*kernel[4]+tmp[8394]*kernel[5]+tmp[8492]*kernel[6]+tmp[8493]*kernel[7]+tmp[8494]*kernel[8];
				ans[8394]<=tmp[8293]*kernel[0]+tmp[8294]*kernel[1]+tmp[8295]*kernel[2]+tmp[8393]*kernel[3]+tmp[8394]*kernel[4]+tmp[8395]*kernel[5]+tmp[8493]*kernel[6]+tmp[8494]*kernel[7]+tmp[8495]*kernel[8];
				ans[8395]<=tmp[8294]*kernel[0]+tmp[8295]*kernel[1]+tmp[8296]*kernel[2]+tmp[8394]*kernel[3]+tmp[8395]*kernel[4]+tmp[8396]*kernel[5]+tmp[8494]*kernel[6]+tmp[8495]*kernel[7]+tmp[8496]*kernel[8];
				ans[8396]<=tmp[8295]*kernel[0]+tmp[8296]*kernel[1]+tmp[8297]*kernel[2]+tmp[8395]*kernel[3]+tmp[8396]*kernel[4]+tmp[8397]*kernel[5]+tmp[8495]*kernel[6]+tmp[8496]*kernel[7]+tmp[8497]*kernel[8];
				ans[8397]<=tmp[8296]*kernel[0]+tmp[8297]*kernel[1]+tmp[8298]*kernel[2]+tmp[8396]*kernel[3]+tmp[8397]*kernel[4]+tmp[8398]*kernel[5]+tmp[8496]*kernel[6]+tmp[8497]*kernel[7]+tmp[8498]*kernel[8];
				ans[8398]<=tmp[8297]*kernel[0]+tmp[8298]*kernel[1]+tmp[8299]*kernel[2]+tmp[8397]*kernel[3]+tmp[8398]*kernel[4]+tmp[8399]*kernel[5]+tmp[8497]*kernel[6]+tmp[8498]*kernel[7]+tmp[8499]*kernel[8];
				ans[8399]<=tmp[8298]*kernel[0]+tmp[8299]*kernel[1]+tmp[8398]*kernel[3]+tmp[8399]*kernel[4]+tmp[8498]*kernel[6]+tmp[8499]*kernel[7];
				ans[8400]<=tmp[8300]*kernel[1]+tmp[8301]*kernel[2]+tmp[8400]*kernel[4]+tmp[8401]*kernel[5]+tmp[8500]*kernel[7]+tmp[8501]*kernel[8];
				ans[8401]<=tmp[8300]*kernel[0]+tmp[8301]*kernel[1]+tmp[8302]*kernel[2]+tmp[8400]*kernel[3]+tmp[8401]*kernel[4]+tmp[8402]*kernel[5]+tmp[8500]*kernel[6]+tmp[8501]*kernel[7]+tmp[8502]*kernel[8];
				ans[8402]<=tmp[8301]*kernel[0]+tmp[8302]*kernel[1]+tmp[8303]*kernel[2]+tmp[8401]*kernel[3]+tmp[8402]*kernel[4]+tmp[8403]*kernel[5]+tmp[8501]*kernel[6]+tmp[8502]*kernel[7]+tmp[8503]*kernel[8];
				ans[8403]<=tmp[8302]*kernel[0]+tmp[8303]*kernel[1]+tmp[8304]*kernel[2]+tmp[8402]*kernel[3]+tmp[8403]*kernel[4]+tmp[8404]*kernel[5]+tmp[8502]*kernel[6]+tmp[8503]*kernel[7]+tmp[8504]*kernel[8];
				ans[8404]<=tmp[8303]*kernel[0]+tmp[8304]*kernel[1]+tmp[8305]*kernel[2]+tmp[8403]*kernel[3]+tmp[8404]*kernel[4]+tmp[8405]*kernel[5]+tmp[8503]*kernel[6]+tmp[8504]*kernel[7]+tmp[8505]*kernel[8];
				ans[8405]<=tmp[8304]*kernel[0]+tmp[8305]*kernel[1]+tmp[8306]*kernel[2]+tmp[8404]*kernel[3]+tmp[8405]*kernel[4]+tmp[8406]*kernel[5]+tmp[8504]*kernel[6]+tmp[8505]*kernel[7]+tmp[8506]*kernel[8];
				ans[8406]<=tmp[8305]*kernel[0]+tmp[8306]*kernel[1]+tmp[8307]*kernel[2]+tmp[8405]*kernel[3]+tmp[8406]*kernel[4]+tmp[8407]*kernel[5]+tmp[8505]*kernel[6]+tmp[8506]*kernel[7]+tmp[8507]*kernel[8];
				ans[8407]<=tmp[8306]*kernel[0]+tmp[8307]*kernel[1]+tmp[8308]*kernel[2]+tmp[8406]*kernel[3]+tmp[8407]*kernel[4]+tmp[8408]*kernel[5]+tmp[8506]*kernel[6]+tmp[8507]*kernel[7]+tmp[8508]*kernel[8];
				ans[8408]<=tmp[8307]*kernel[0]+tmp[8308]*kernel[1]+tmp[8309]*kernel[2]+tmp[8407]*kernel[3]+tmp[8408]*kernel[4]+tmp[8409]*kernel[5]+tmp[8507]*kernel[6]+tmp[8508]*kernel[7]+tmp[8509]*kernel[8];
				ans[8409]<=tmp[8308]*kernel[0]+tmp[8309]*kernel[1]+tmp[8310]*kernel[2]+tmp[8408]*kernel[3]+tmp[8409]*kernel[4]+tmp[8410]*kernel[5]+tmp[8508]*kernel[6]+tmp[8509]*kernel[7]+tmp[8510]*kernel[8];
				ans[8410]<=tmp[8309]*kernel[0]+tmp[8310]*kernel[1]+tmp[8311]*kernel[2]+tmp[8409]*kernel[3]+tmp[8410]*kernel[4]+tmp[8411]*kernel[5]+tmp[8509]*kernel[6]+tmp[8510]*kernel[7]+tmp[8511]*kernel[8];
				ans[8411]<=tmp[8310]*kernel[0]+tmp[8311]*kernel[1]+tmp[8312]*kernel[2]+tmp[8410]*kernel[3]+tmp[8411]*kernel[4]+tmp[8412]*kernel[5]+tmp[8510]*kernel[6]+tmp[8511]*kernel[7]+tmp[8512]*kernel[8];
				ans[8412]<=tmp[8311]*kernel[0]+tmp[8312]*kernel[1]+tmp[8313]*kernel[2]+tmp[8411]*kernel[3]+tmp[8412]*kernel[4]+tmp[8413]*kernel[5]+tmp[8511]*kernel[6]+tmp[8512]*kernel[7]+tmp[8513]*kernel[8];
				ans[8413]<=tmp[8312]*kernel[0]+tmp[8313]*kernel[1]+tmp[8314]*kernel[2]+tmp[8412]*kernel[3]+tmp[8413]*kernel[4]+tmp[8414]*kernel[5]+tmp[8512]*kernel[6]+tmp[8513]*kernel[7]+tmp[8514]*kernel[8];
				ans[8414]<=tmp[8313]*kernel[0]+tmp[8314]*kernel[1]+tmp[8315]*kernel[2]+tmp[8413]*kernel[3]+tmp[8414]*kernel[4]+tmp[8415]*kernel[5]+tmp[8513]*kernel[6]+tmp[8514]*kernel[7]+tmp[8515]*kernel[8];
				ans[8415]<=tmp[8314]*kernel[0]+tmp[8315]*kernel[1]+tmp[8316]*kernel[2]+tmp[8414]*kernel[3]+tmp[8415]*kernel[4]+tmp[8416]*kernel[5]+tmp[8514]*kernel[6]+tmp[8515]*kernel[7]+tmp[8516]*kernel[8];
				ans[8416]<=tmp[8315]*kernel[0]+tmp[8316]*kernel[1]+tmp[8317]*kernel[2]+tmp[8415]*kernel[3]+tmp[8416]*kernel[4]+tmp[8417]*kernel[5]+tmp[8515]*kernel[6]+tmp[8516]*kernel[7]+tmp[8517]*kernel[8];
				ans[8417]<=tmp[8316]*kernel[0]+tmp[8317]*kernel[1]+tmp[8318]*kernel[2]+tmp[8416]*kernel[3]+tmp[8417]*kernel[4]+tmp[8418]*kernel[5]+tmp[8516]*kernel[6]+tmp[8517]*kernel[7]+tmp[8518]*kernel[8];
				ans[8418]<=tmp[8317]*kernel[0]+tmp[8318]*kernel[1]+tmp[8319]*kernel[2]+tmp[8417]*kernel[3]+tmp[8418]*kernel[4]+tmp[8419]*kernel[5]+tmp[8517]*kernel[6]+tmp[8518]*kernel[7]+tmp[8519]*kernel[8];
				ans[8419]<=tmp[8318]*kernel[0]+tmp[8319]*kernel[1]+tmp[8320]*kernel[2]+tmp[8418]*kernel[3]+tmp[8419]*kernel[4]+tmp[8420]*kernel[5]+tmp[8518]*kernel[6]+tmp[8519]*kernel[7]+tmp[8520]*kernel[8];
				ans[8420]<=tmp[8319]*kernel[0]+tmp[8320]*kernel[1]+tmp[8321]*kernel[2]+tmp[8419]*kernel[3]+tmp[8420]*kernel[4]+tmp[8421]*kernel[5]+tmp[8519]*kernel[6]+tmp[8520]*kernel[7]+tmp[8521]*kernel[8];
				ans[8421]<=tmp[8320]*kernel[0]+tmp[8321]*kernel[1]+tmp[8322]*kernel[2]+tmp[8420]*kernel[3]+tmp[8421]*kernel[4]+tmp[8422]*kernel[5]+tmp[8520]*kernel[6]+tmp[8521]*kernel[7]+tmp[8522]*kernel[8];
				ans[8422]<=tmp[8321]*kernel[0]+tmp[8322]*kernel[1]+tmp[8323]*kernel[2]+tmp[8421]*kernel[3]+tmp[8422]*kernel[4]+tmp[8423]*kernel[5]+tmp[8521]*kernel[6]+tmp[8522]*kernel[7]+tmp[8523]*kernel[8];
				ans[8423]<=tmp[8322]*kernel[0]+tmp[8323]*kernel[1]+tmp[8324]*kernel[2]+tmp[8422]*kernel[3]+tmp[8423]*kernel[4]+tmp[8424]*kernel[5]+tmp[8522]*kernel[6]+tmp[8523]*kernel[7]+tmp[8524]*kernel[8];
				ans[8424]<=tmp[8323]*kernel[0]+tmp[8324]*kernel[1]+tmp[8325]*kernel[2]+tmp[8423]*kernel[3]+tmp[8424]*kernel[4]+tmp[8425]*kernel[5]+tmp[8523]*kernel[6]+tmp[8524]*kernel[7]+tmp[8525]*kernel[8];
				ans[8425]<=tmp[8324]*kernel[0]+tmp[8325]*kernel[1]+tmp[8326]*kernel[2]+tmp[8424]*kernel[3]+tmp[8425]*kernel[4]+tmp[8426]*kernel[5]+tmp[8524]*kernel[6]+tmp[8525]*kernel[7]+tmp[8526]*kernel[8];
				ans[8426]<=tmp[8325]*kernel[0]+tmp[8326]*kernel[1]+tmp[8327]*kernel[2]+tmp[8425]*kernel[3]+tmp[8426]*kernel[4]+tmp[8427]*kernel[5]+tmp[8525]*kernel[6]+tmp[8526]*kernel[7]+tmp[8527]*kernel[8];
				ans[8427]<=tmp[8326]*kernel[0]+tmp[8327]*kernel[1]+tmp[8328]*kernel[2]+tmp[8426]*kernel[3]+tmp[8427]*kernel[4]+tmp[8428]*kernel[5]+tmp[8526]*kernel[6]+tmp[8527]*kernel[7]+tmp[8528]*kernel[8];
				ans[8428]<=tmp[8327]*kernel[0]+tmp[8328]*kernel[1]+tmp[8329]*kernel[2]+tmp[8427]*kernel[3]+tmp[8428]*kernel[4]+tmp[8429]*kernel[5]+tmp[8527]*kernel[6]+tmp[8528]*kernel[7]+tmp[8529]*kernel[8];
				ans[8429]<=tmp[8328]*kernel[0]+tmp[8329]*kernel[1]+tmp[8330]*kernel[2]+tmp[8428]*kernel[3]+tmp[8429]*kernel[4]+tmp[8430]*kernel[5]+tmp[8528]*kernel[6]+tmp[8529]*kernel[7]+tmp[8530]*kernel[8];
				ans[8430]<=tmp[8329]*kernel[0]+tmp[8330]*kernel[1]+tmp[8331]*kernel[2]+tmp[8429]*kernel[3]+tmp[8430]*kernel[4]+tmp[8431]*kernel[5]+tmp[8529]*kernel[6]+tmp[8530]*kernel[7]+tmp[8531]*kernel[8];
				ans[8431]<=tmp[8330]*kernel[0]+tmp[8331]*kernel[1]+tmp[8332]*kernel[2]+tmp[8430]*kernel[3]+tmp[8431]*kernel[4]+tmp[8432]*kernel[5]+tmp[8530]*kernel[6]+tmp[8531]*kernel[7]+tmp[8532]*kernel[8];
				ans[8432]<=tmp[8331]*kernel[0]+tmp[8332]*kernel[1]+tmp[8333]*kernel[2]+tmp[8431]*kernel[3]+tmp[8432]*kernel[4]+tmp[8433]*kernel[5]+tmp[8531]*kernel[6]+tmp[8532]*kernel[7]+tmp[8533]*kernel[8];
				ans[8433]<=tmp[8332]*kernel[0]+tmp[8333]*kernel[1]+tmp[8334]*kernel[2]+tmp[8432]*kernel[3]+tmp[8433]*kernel[4]+tmp[8434]*kernel[5]+tmp[8532]*kernel[6]+tmp[8533]*kernel[7]+tmp[8534]*kernel[8];
				ans[8434]<=tmp[8333]*kernel[0]+tmp[8334]*kernel[1]+tmp[8335]*kernel[2]+tmp[8433]*kernel[3]+tmp[8434]*kernel[4]+tmp[8435]*kernel[5]+tmp[8533]*kernel[6]+tmp[8534]*kernel[7]+tmp[8535]*kernel[8];
				ans[8435]<=tmp[8334]*kernel[0]+tmp[8335]*kernel[1]+tmp[8336]*kernel[2]+tmp[8434]*kernel[3]+tmp[8435]*kernel[4]+tmp[8436]*kernel[5]+tmp[8534]*kernel[6]+tmp[8535]*kernel[7]+tmp[8536]*kernel[8];
				ans[8436]<=tmp[8335]*kernel[0]+tmp[8336]*kernel[1]+tmp[8337]*kernel[2]+tmp[8435]*kernel[3]+tmp[8436]*kernel[4]+tmp[8437]*kernel[5]+tmp[8535]*kernel[6]+tmp[8536]*kernel[7]+tmp[8537]*kernel[8];
				ans[8437]<=tmp[8336]*kernel[0]+tmp[8337]*kernel[1]+tmp[8338]*kernel[2]+tmp[8436]*kernel[3]+tmp[8437]*kernel[4]+tmp[8438]*kernel[5]+tmp[8536]*kernel[6]+tmp[8537]*kernel[7]+tmp[8538]*kernel[8];
				ans[8438]<=tmp[8337]*kernel[0]+tmp[8338]*kernel[1]+tmp[8339]*kernel[2]+tmp[8437]*kernel[3]+tmp[8438]*kernel[4]+tmp[8439]*kernel[5]+tmp[8537]*kernel[6]+tmp[8538]*kernel[7]+tmp[8539]*kernel[8];
				ans[8439]<=tmp[8338]*kernel[0]+tmp[8339]*kernel[1]+tmp[8340]*kernel[2]+tmp[8438]*kernel[3]+tmp[8439]*kernel[4]+tmp[8440]*kernel[5]+tmp[8538]*kernel[6]+tmp[8539]*kernel[7]+tmp[8540]*kernel[8];
				ans[8440]<=tmp[8339]*kernel[0]+tmp[8340]*kernel[1]+tmp[8341]*kernel[2]+tmp[8439]*kernel[3]+tmp[8440]*kernel[4]+tmp[8441]*kernel[5]+tmp[8539]*kernel[6]+tmp[8540]*kernel[7]+tmp[8541]*kernel[8];
				ans[8441]<=tmp[8340]*kernel[0]+tmp[8341]*kernel[1]+tmp[8342]*kernel[2]+tmp[8440]*kernel[3]+tmp[8441]*kernel[4]+tmp[8442]*kernel[5]+tmp[8540]*kernel[6]+tmp[8541]*kernel[7]+tmp[8542]*kernel[8];
				ans[8442]<=tmp[8341]*kernel[0]+tmp[8342]*kernel[1]+tmp[8343]*kernel[2]+tmp[8441]*kernel[3]+tmp[8442]*kernel[4]+tmp[8443]*kernel[5]+tmp[8541]*kernel[6]+tmp[8542]*kernel[7]+tmp[8543]*kernel[8];
				ans[8443]<=tmp[8342]*kernel[0]+tmp[8343]*kernel[1]+tmp[8344]*kernel[2]+tmp[8442]*kernel[3]+tmp[8443]*kernel[4]+tmp[8444]*kernel[5]+tmp[8542]*kernel[6]+tmp[8543]*kernel[7]+tmp[8544]*kernel[8];
				ans[8444]<=tmp[8343]*kernel[0]+tmp[8344]*kernel[1]+tmp[8345]*kernel[2]+tmp[8443]*kernel[3]+tmp[8444]*kernel[4]+tmp[8445]*kernel[5]+tmp[8543]*kernel[6]+tmp[8544]*kernel[7]+tmp[8545]*kernel[8];
				ans[8445]<=tmp[8344]*kernel[0]+tmp[8345]*kernel[1]+tmp[8346]*kernel[2]+tmp[8444]*kernel[3]+tmp[8445]*kernel[4]+tmp[8446]*kernel[5]+tmp[8544]*kernel[6]+tmp[8545]*kernel[7]+tmp[8546]*kernel[8];
				ans[8446]<=tmp[8345]*kernel[0]+tmp[8346]*kernel[1]+tmp[8347]*kernel[2]+tmp[8445]*kernel[3]+tmp[8446]*kernel[4]+tmp[8447]*kernel[5]+tmp[8545]*kernel[6]+tmp[8546]*kernel[7]+tmp[8547]*kernel[8];
				ans[8447]<=tmp[8346]*kernel[0]+tmp[8347]*kernel[1]+tmp[8348]*kernel[2]+tmp[8446]*kernel[3]+tmp[8447]*kernel[4]+tmp[8448]*kernel[5]+tmp[8546]*kernel[6]+tmp[8547]*kernel[7]+tmp[8548]*kernel[8];
				ans[8448]<=tmp[8347]*kernel[0]+tmp[8348]*kernel[1]+tmp[8349]*kernel[2]+tmp[8447]*kernel[3]+tmp[8448]*kernel[4]+tmp[8449]*kernel[5]+tmp[8547]*kernel[6]+tmp[8548]*kernel[7]+tmp[8549]*kernel[8];
				ans[8449]<=tmp[8348]*kernel[0]+tmp[8349]*kernel[1]+tmp[8350]*kernel[2]+tmp[8448]*kernel[3]+tmp[8449]*kernel[4]+tmp[8450]*kernel[5]+tmp[8548]*kernel[6]+tmp[8549]*kernel[7]+tmp[8550]*kernel[8];
				ans[8450]<=tmp[8349]*kernel[0]+tmp[8350]*kernel[1]+tmp[8351]*kernel[2]+tmp[8449]*kernel[3]+tmp[8450]*kernel[4]+tmp[8451]*kernel[5]+tmp[8549]*kernel[6]+tmp[8550]*kernel[7]+tmp[8551]*kernel[8];
				ans[8451]<=tmp[8350]*kernel[0]+tmp[8351]*kernel[1]+tmp[8352]*kernel[2]+tmp[8450]*kernel[3]+tmp[8451]*kernel[4]+tmp[8452]*kernel[5]+tmp[8550]*kernel[6]+tmp[8551]*kernel[7]+tmp[8552]*kernel[8];
				ans[8452]<=tmp[8351]*kernel[0]+tmp[8352]*kernel[1]+tmp[8353]*kernel[2]+tmp[8451]*kernel[3]+tmp[8452]*kernel[4]+tmp[8453]*kernel[5]+tmp[8551]*kernel[6]+tmp[8552]*kernel[7]+tmp[8553]*kernel[8];
				ans[8453]<=tmp[8352]*kernel[0]+tmp[8353]*kernel[1]+tmp[8354]*kernel[2]+tmp[8452]*kernel[3]+tmp[8453]*kernel[4]+tmp[8454]*kernel[5]+tmp[8552]*kernel[6]+tmp[8553]*kernel[7]+tmp[8554]*kernel[8];
				ans[8454]<=tmp[8353]*kernel[0]+tmp[8354]*kernel[1]+tmp[8355]*kernel[2]+tmp[8453]*kernel[3]+tmp[8454]*kernel[4]+tmp[8455]*kernel[5]+tmp[8553]*kernel[6]+tmp[8554]*kernel[7]+tmp[8555]*kernel[8];
				ans[8455]<=tmp[8354]*kernel[0]+tmp[8355]*kernel[1]+tmp[8356]*kernel[2]+tmp[8454]*kernel[3]+tmp[8455]*kernel[4]+tmp[8456]*kernel[5]+tmp[8554]*kernel[6]+tmp[8555]*kernel[7]+tmp[8556]*kernel[8];
				ans[8456]<=tmp[8355]*kernel[0]+tmp[8356]*kernel[1]+tmp[8357]*kernel[2]+tmp[8455]*kernel[3]+tmp[8456]*kernel[4]+tmp[8457]*kernel[5]+tmp[8555]*kernel[6]+tmp[8556]*kernel[7]+tmp[8557]*kernel[8];
				ans[8457]<=tmp[8356]*kernel[0]+tmp[8357]*kernel[1]+tmp[8358]*kernel[2]+tmp[8456]*kernel[3]+tmp[8457]*kernel[4]+tmp[8458]*kernel[5]+tmp[8556]*kernel[6]+tmp[8557]*kernel[7]+tmp[8558]*kernel[8];
				ans[8458]<=tmp[8357]*kernel[0]+tmp[8358]*kernel[1]+tmp[8359]*kernel[2]+tmp[8457]*kernel[3]+tmp[8458]*kernel[4]+tmp[8459]*kernel[5]+tmp[8557]*kernel[6]+tmp[8558]*kernel[7]+tmp[8559]*kernel[8];
				ans[8459]<=tmp[8358]*kernel[0]+tmp[8359]*kernel[1]+tmp[8360]*kernel[2]+tmp[8458]*kernel[3]+tmp[8459]*kernel[4]+tmp[8460]*kernel[5]+tmp[8558]*kernel[6]+tmp[8559]*kernel[7]+tmp[8560]*kernel[8];
				ans[8460]<=tmp[8359]*kernel[0]+tmp[8360]*kernel[1]+tmp[8361]*kernel[2]+tmp[8459]*kernel[3]+tmp[8460]*kernel[4]+tmp[8461]*kernel[5]+tmp[8559]*kernel[6]+tmp[8560]*kernel[7]+tmp[8561]*kernel[8];
				ans[8461]<=tmp[8360]*kernel[0]+tmp[8361]*kernel[1]+tmp[8362]*kernel[2]+tmp[8460]*kernel[3]+tmp[8461]*kernel[4]+tmp[8462]*kernel[5]+tmp[8560]*kernel[6]+tmp[8561]*kernel[7]+tmp[8562]*kernel[8];
				ans[8462]<=tmp[8361]*kernel[0]+tmp[8362]*kernel[1]+tmp[8363]*kernel[2]+tmp[8461]*kernel[3]+tmp[8462]*kernel[4]+tmp[8463]*kernel[5]+tmp[8561]*kernel[6]+tmp[8562]*kernel[7]+tmp[8563]*kernel[8];
				ans[8463]<=tmp[8362]*kernel[0]+tmp[8363]*kernel[1]+tmp[8364]*kernel[2]+tmp[8462]*kernel[3]+tmp[8463]*kernel[4]+tmp[8464]*kernel[5]+tmp[8562]*kernel[6]+tmp[8563]*kernel[7]+tmp[8564]*kernel[8];
				ans[8464]<=tmp[8363]*kernel[0]+tmp[8364]*kernel[1]+tmp[8365]*kernel[2]+tmp[8463]*kernel[3]+tmp[8464]*kernel[4]+tmp[8465]*kernel[5]+tmp[8563]*kernel[6]+tmp[8564]*kernel[7]+tmp[8565]*kernel[8];
				ans[8465]<=tmp[8364]*kernel[0]+tmp[8365]*kernel[1]+tmp[8366]*kernel[2]+tmp[8464]*kernel[3]+tmp[8465]*kernel[4]+tmp[8466]*kernel[5]+tmp[8564]*kernel[6]+tmp[8565]*kernel[7]+tmp[8566]*kernel[8];
				ans[8466]<=tmp[8365]*kernel[0]+tmp[8366]*kernel[1]+tmp[8367]*kernel[2]+tmp[8465]*kernel[3]+tmp[8466]*kernel[4]+tmp[8467]*kernel[5]+tmp[8565]*kernel[6]+tmp[8566]*kernel[7]+tmp[8567]*kernel[8];
				ans[8467]<=tmp[8366]*kernel[0]+tmp[8367]*kernel[1]+tmp[8368]*kernel[2]+tmp[8466]*kernel[3]+tmp[8467]*kernel[4]+tmp[8468]*kernel[5]+tmp[8566]*kernel[6]+tmp[8567]*kernel[7]+tmp[8568]*kernel[8];
				ans[8468]<=tmp[8367]*kernel[0]+tmp[8368]*kernel[1]+tmp[8369]*kernel[2]+tmp[8467]*kernel[3]+tmp[8468]*kernel[4]+tmp[8469]*kernel[5]+tmp[8567]*kernel[6]+tmp[8568]*kernel[7]+tmp[8569]*kernel[8];
				ans[8469]<=tmp[8368]*kernel[0]+tmp[8369]*kernel[1]+tmp[8370]*kernel[2]+tmp[8468]*kernel[3]+tmp[8469]*kernel[4]+tmp[8470]*kernel[5]+tmp[8568]*kernel[6]+tmp[8569]*kernel[7]+tmp[8570]*kernel[8];
				ans[8470]<=tmp[8369]*kernel[0]+tmp[8370]*kernel[1]+tmp[8371]*kernel[2]+tmp[8469]*kernel[3]+tmp[8470]*kernel[4]+tmp[8471]*kernel[5]+tmp[8569]*kernel[6]+tmp[8570]*kernel[7]+tmp[8571]*kernel[8];
				ans[8471]<=tmp[8370]*kernel[0]+tmp[8371]*kernel[1]+tmp[8372]*kernel[2]+tmp[8470]*kernel[3]+tmp[8471]*kernel[4]+tmp[8472]*kernel[5]+tmp[8570]*kernel[6]+tmp[8571]*kernel[7]+tmp[8572]*kernel[8];
				ans[8472]<=tmp[8371]*kernel[0]+tmp[8372]*kernel[1]+tmp[8373]*kernel[2]+tmp[8471]*kernel[3]+tmp[8472]*kernel[4]+tmp[8473]*kernel[5]+tmp[8571]*kernel[6]+tmp[8572]*kernel[7]+tmp[8573]*kernel[8];
				ans[8473]<=tmp[8372]*kernel[0]+tmp[8373]*kernel[1]+tmp[8374]*kernel[2]+tmp[8472]*kernel[3]+tmp[8473]*kernel[4]+tmp[8474]*kernel[5]+tmp[8572]*kernel[6]+tmp[8573]*kernel[7]+tmp[8574]*kernel[8];
				ans[8474]<=tmp[8373]*kernel[0]+tmp[8374]*kernel[1]+tmp[8375]*kernel[2]+tmp[8473]*kernel[3]+tmp[8474]*kernel[4]+tmp[8475]*kernel[5]+tmp[8573]*kernel[6]+tmp[8574]*kernel[7]+tmp[8575]*kernel[8];
				ans[8475]<=tmp[8374]*kernel[0]+tmp[8375]*kernel[1]+tmp[8376]*kernel[2]+tmp[8474]*kernel[3]+tmp[8475]*kernel[4]+tmp[8476]*kernel[5]+tmp[8574]*kernel[6]+tmp[8575]*kernel[7]+tmp[8576]*kernel[8];
				ans[8476]<=tmp[8375]*kernel[0]+tmp[8376]*kernel[1]+tmp[8377]*kernel[2]+tmp[8475]*kernel[3]+tmp[8476]*kernel[4]+tmp[8477]*kernel[5]+tmp[8575]*kernel[6]+tmp[8576]*kernel[7]+tmp[8577]*kernel[8];
				ans[8477]<=tmp[8376]*kernel[0]+tmp[8377]*kernel[1]+tmp[8378]*kernel[2]+tmp[8476]*kernel[3]+tmp[8477]*kernel[4]+tmp[8478]*kernel[5]+tmp[8576]*kernel[6]+tmp[8577]*kernel[7]+tmp[8578]*kernel[8];
				ans[8478]<=tmp[8377]*kernel[0]+tmp[8378]*kernel[1]+tmp[8379]*kernel[2]+tmp[8477]*kernel[3]+tmp[8478]*kernel[4]+tmp[8479]*kernel[5]+tmp[8577]*kernel[6]+tmp[8578]*kernel[7]+tmp[8579]*kernel[8];
				ans[8479]<=tmp[8378]*kernel[0]+tmp[8379]*kernel[1]+tmp[8380]*kernel[2]+tmp[8478]*kernel[3]+tmp[8479]*kernel[4]+tmp[8480]*kernel[5]+tmp[8578]*kernel[6]+tmp[8579]*kernel[7]+tmp[8580]*kernel[8];
				ans[8480]<=tmp[8379]*kernel[0]+tmp[8380]*kernel[1]+tmp[8381]*kernel[2]+tmp[8479]*kernel[3]+tmp[8480]*kernel[4]+tmp[8481]*kernel[5]+tmp[8579]*kernel[6]+tmp[8580]*kernel[7]+tmp[8581]*kernel[8];
				ans[8481]<=tmp[8380]*kernel[0]+tmp[8381]*kernel[1]+tmp[8382]*kernel[2]+tmp[8480]*kernel[3]+tmp[8481]*kernel[4]+tmp[8482]*kernel[5]+tmp[8580]*kernel[6]+tmp[8581]*kernel[7]+tmp[8582]*kernel[8];
				ans[8482]<=tmp[8381]*kernel[0]+tmp[8382]*kernel[1]+tmp[8383]*kernel[2]+tmp[8481]*kernel[3]+tmp[8482]*kernel[4]+tmp[8483]*kernel[5]+tmp[8581]*kernel[6]+tmp[8582]*kernel[7]+tmp[8583]*kernel[8];
				ans[8483]<=tmp[8382]*kernel[0]+tmp[8383]*kernel[1]+tmp[8384]*kernel[2]+tmp[8482]*kernel[3]+tmp[8483]*kernel[4]+tmp[8484]*kernel[5]+tmp[8582]*kernel[6]+tmp[8583]*kernel[7]+tmp[8584]*kernel[8];
				ans[8484]<=tmp[8383]*kernel[0]+tmp[8384]*kernel[1]+tmp[8385]*kernel[2]+tmp[8483]*kernel[3]+tmp[8484]*kernel[4]+tmp[8485]*kernel[5]+tmp[8583]*kernel[6]+tmp[8584]*kernel[7]+tmp[8585]*kernel[8];
				ans[8485]<=tmp[8384]*kernel[0]+tmp[8385]*kernel[1]+tmp[8386]*kernel[2]+tmp[8484]*kernel[3]+tmp[8485]*kernel[4]+tmp[8486]*kernel[5]+tmp[8584]*kernel[6]+tmp[8585]*kernel[7]+tmp[8586]*kernel[8];
				ans[8486]<=tmp[8385]*kernel[0]+tmp[8386]*kernel[1]+tmp[8387]*kernel[2]+tmp[8485]*kernel[3]+tmp[8486]*kernel[4]+tmp[8487]*kernel[5]+tmp[8585]*kernel[6]+tmp[8586]*kernel[7]+tmp[8587]*kernel[8];
				ans[8487]<=tmp[8386]*kernel[0]+tmp[8387]*kernel[1]+tmp[8388]*kernel[2]+tmp[8486]*kernel[3]+tmp[8487]*kernel[4]+tmp[8488]*kernel[5]+tmp[8586]*kernel[6]+tmp[8587]*kernel[7]+tmp[8588]*kernel[8];
				ans[8488]<=tmp[8387]*kernel[0]+tmp[8388]*kernel[1]+tmp[8389]*kernel[2]+tmp[8487]*kernel[3]+tmp[8488]*kernel[4]+tmp[8489]*kernel[5]+tmp[8587]*kernel[6]+tmp[8588]*kernel[7]+tmp[8589]*kernel[8];
				ans[8489]<=tmp[8388]*kernel[0]+tmp[8389]*kernel[1]+tmp[8390]*kernel[2]+tmp[8488]*kernel[3]+tmp[8489]*kernel[4]+tmp[8490]*kernel[5]+tmp[8588]*kernel[6]+tmp[8589]*kernel[7]+tmp[8590]*kernel[8];
				ans[8490]<=tmp[8389]*kernel[0]+tmp[8390]*kernel[1]+tmp[8391]*kernel[2]+tmp[8489]*kernel[3]+tmp[8490]*kernel[4]+tmp[8491]*kernel[5]+tmp[8589]*kernel[6]+tmp[8590]*kernel[7]+tmp[8591]*kernel[8];
				ans[8491]<=tmp[8390]*kernel[0]+tmp[8391]*kernel[1]+tmp[8392]*kernel[2]+tmp[8490]*kernel[3]+tmp[8491]*kernel[4]+tmp[8492]*kernel[5]+tmp[8590]*kernel[6]+tmp[8591]*kernel[7]+tmp[8592]*kernel[8];
				ans[8492]<=tmp[8391]*kernel[0]+tmp[8392]*kernel[1]+tmp[8393]*kernel[2]+tmp[8491]*kernel[3]+tmp[8492]*kernel[4]+tmp[8493]*kernel[5]+tmp[8591]*kernel[6]+tmp[8592]*kernel[7]+tmp[8593]*kernel[8];
				ans[8493]<=tmp[8392]*kernel[0]+tmp[8393]*kernel[1]+tmp[8394]*kernel[2]+tmp[8492]*kernel[3]+tmp[8493]*kernel[4]+tmp[8494]*kernel[5]+tmp[8592]*kernel[6]+tmp[8593]*kernel[7]+tmp[8594]*kernel[8];
				ans[8494]<=tmp[8393]*kernel[0]+tmp[8394]*kernel[1]+tmp[8395]*kernel[2]+tmp[8493]*kernel[3]+tmp[8494]*kernel[4]+tmp[8495]*kernel[5]+tmp[8593]*kernel[6]+tmp[8594]*kernel[7]+tmp[8595]*kernel[8];
				ans[8495]<=tmp[8394]*kernel[0]+tmp[8395]*kernel[1]+tmp[8396]*kernel[2]+tmp[8494]*kernel[3]+tmp[8495]*kernel[4]+tmp[8496]*kernel[5]+tmp[8594]*kernel[6]+tmp[8595]*kernel[7]+tmp[8596]*kernel[8];
				ans[8496]<=tmp[8395]*kernel[0]+tmp[8396]*kernel[1]+tmp[8397]*kernel[2]+tmp[8495]*kernel[3]+tmp[8496]*kernel[4]+tmp[8497]*kernel[5]+tmp[8595]*kernel[6]+tmp[8596]*kernel[7]+tmp[8597]*kernel[8];
				ans[8497]<=tmp[8396]*kernel[0]+tmp[8397]*kernel[1]+tmp[8398]*kernel[2]+tmp[8496]*kernel[3]+tmp[8497]*kernel[4]+tmp[8498]*kernel[5]+tmp[8596]*kernel[6]+tmp[8597]*kernel[7]+tmp[8598]*kernel[8];
				ans[8498]<=tmp[8397]*kernel[0]+tmp[8398]*kernel[1]+tmp[8399]*kernel[2]+tmp[8497]*kernel[3]+tmp[8498]*kernel[4]+tmp[8499]*kernel[5]+tmp[8597]*kernel[6]+tmp[8598]*kernel[7]+tmp[8599]*kernel[8];
				ans[8499]<=tmp[8398]*kernel[0]+tmp[8399]*kernel[1]+tmp[8498]*kernel[3]+tmp[8499]*kernel[4]+tmp[8598]*kernel[6]+tmp[8599]*kernel[7];
				ans[8500]<=tmp[8400]*kernel[1]+tmp[8401]*kernel[2]+tmp[8500]*kernel[4]+tmp[8501]*kernel[5]+tmp[8600]*kernel[7]+tmp[8601]*kernel[8];
				ans[8501]<=tmp[8400]*kernel[0]+tmp[8401]*kernel[1]+tmp[8402]*kernel[2]+tmp[8500]*kernel[3]+tmp[8501]*kernel[4]+tmp[8502]*kernel[5]+tmp[8600]*kernel[6]+tmp[8601]*kernel[7]+tmp[8602]*kernel[8];
				ans[8502]<=tmp[8401]*kernel[0]+tmp[8402]*kernel[1]+tmp[8403]*kernel[2]+tmp[8501]*kernel[3]+tmp[8502]*kernel[4]+tmp[8503]*kernel[5]+tmp[8601]*kernel[6]+tmp[8602]*kernel[7]+tmp[8603]*kernel[8];
				ans[8503]<=tmp[8402]*kernel[0]+tmp[8403]*kernel[1]+tmp[8404]*kernel[2]+tmp[8502]*kernel[3]+tmp[8503]*kernel[4]+tmp[8504]*kernel[5]+tmp[8602]*kernel[6]+tmp[8603]*kernel[7]+tmp[8604]*kernel[8];
				ans[8504]<=tmp[8403]*kernel[0]+tmp[8404]*kernel[1]+tmp[8405]*kernel[2]+tmp[8503]*kernel[3]+tmp[8504]*kernel[4]+tmp[8505]*kernel[5]+tmp[8603]*kernel[6]+tmp[8604]*kernel[7]+tmp[8605]*kernel[8];
				ans[8505]<=tmp[8404]*kernel[0]+tmp[8405]*kernel[1]+tmp[8406]*kernel[2]+tmp[8504]*kernel[3]+tmp[8505]*kernel[4]+tmp[8506]*kernel[5]+tmp[8604]*kernel[6]+tmp[8605]*kernel[7]+tmp[8606]*kernel[8];
				ans[8506]<=tmp[8405]*kernel[0]+tmp[8406]*kernel[1]+tmp[8407]*kernel[2]+tmp[8505]*kernel[3]+tmp[8506]*kernel[4]+tmp[8507]*kernel[5]+tmp[8605]*kernel[6]+tmp[8606]*kernel[7]+tmp[8607]*kernel[8];
				ans[8507]<=tmp[8406]*kernel[0]+tmp[8407]*kernel[1]+tmp[8408]*kernel[2]+tmp[8506]*kernel[3]+tmp[8507]*kernel[4]+tmp[8508]*kernel[5]+tmp[8606]*kernel[6]+tmp[8607]*kernel[7]+tmp[8608]*kernel[8];
				ans[8508]<=tmp[8407]*kernel[0]+tmp[8408]*kernel[1]+tmp[8409]*kernel[2]+tmp[8507]*kernel[3]+tmp[8508]*kernel[4]+tmp[8509]*kernel[5]+tmp[8607]*kernel[6]+tmp[8608]*kernel[7]+tmp[8609]*kernel[8];
				ans[8509]<=tmp[8408]*kernel[0]+tmp[8409]*kernel[1]+tmp[8410]*kernel[2]+tmp[8508]*kernel[3]+tmp[8509]*kernel[4]+tmp[8510]*kernel[5]+tmp[8608]*kernel[6]+tmp[8609]*kernel[7]+tmp[8610]*kernel[8];
				ans[8510]<=tmp[8409]*kernel[0]+tmp[8410]*kernel[1]+tmp[8411]*kernel[2]+tmp[8509]*kernel[3]+tmp[8510]*kernel[4]+tmp[8511]*kernel[5]+tmp[8609]*kernel[6]+tmp[8610]*kernel[7]+tmp[8611]*kernel[8];
				ans[8511]<=tmp[8410]*kernel[0]+tmp[8411]*kernel[1]+tmp[8412]*kernel[2]+tmp[8510]*kernel[3]+tmp[8511]*kernel[4]+tmp[8512]*kernel[5]+tmp[8610]*kernel[6]+tmp[8611]*kernel[7]+tmp[8612]*kernel[8];
				ans[8512]<=tmp[8411]*kernel[0]+tmp[8412]*kernel[1]+tmp[8413]*kernel[2]+tmp[8511]*kernel[3]+tmp[8512]*kernel[4]+tmp[8513]*kernel[5]+tmp[8611]*kernel[6]+tmp[8612]*kernel[7]+tmp[8613]*kernel[8];
				ans[8513]<=tmp[8412]*kernel[0]+tmp[8413]*kernel[1]+tmp[8414]*kernel[2]+tmp[8512]*kernel[3]+tmp[8513]*kernel[4]+tmp[8514]*kernel[5]+tmp[8612]*kernel[6]+tmp[8613]*kernel[7]+tmp[8614]*kernel[8];
				ans[8514]<=tmp[8413]*kernel[0]+tmp[8414]*kernel[1]+tmp[8415]*kernel[2]+tmp[8513]*kernel[3]+tmp[8514]*kernel[4]+tmp[8515]*kernel[5]+tmp[8613]*kernel[6]+tmp[8614]*kernel[7]+tmp[8615]*kernel[8];
				ans[8515]<=tmp[8414]*kernel[0]+tmp[8415]*kernel[1]+tmp[8416]*kernel[2]+tmp[8514]*kernel[3]+tmp[8515]*kernel[4]+tmp[8516]*kernel[5]+tmp[8614]*kernel[6]+tmp[8615]*kernel[7]+tmp[8616]*kernel[8];
				ans[8516]<=tmp[8415]*kernel[0]+tmp[8416]*kernel[1]+tmp[8417]*kernel[2]+tmp[8515]*kernel[3]+tmp[8516]*kernel[4]+tmp[8517]*kernel[5]+tmp[8615]*kernel[6]+tmp[8616]*kernel[7]+tmp[8617]*kernel[8];
				ans[8517]<=tmp[8416]*kernel[0]+tmp[8417]*kernel[1]+tmp[8418]*kernel[2]+tmp[8516]*kernel[3]+tmp[8517]*kernel[4]+tmp[8518]*kernel[5]+tmp[8616]*kernel[6]+tmp[8617]*kernel[7]+tmp[8618]*kernel[8];
				ans[8518]<=tmp[8417]*kernel[0]+tmp[8418]*kernel[1]+tmp[8419]*kernel[2]+tmp[8517]*kernel[3]+tmp[8518]*kernel[4]+tmp[8519]*kernel[5]+tmp[8617]*kernel[6]+tmp[8618]*kernel[7]+tmp[8619]*kernel[8];
				ans[8519]<=tmp[8418]*kernel[0]+tmp[8419]*kernel[1]+tmp[8420]*kernel[2]+tmp[8518]*kernel[3]+tmp[8519]*kernel[4]+tmp[8520]*kernel[5]+tmp[8618]*kernel[6]+tmp[8619]*kernel[7]+tmp[8620]*kernel[8];
				ans[8520]<=tmp[8419]*kernel[0]+tmp[8420]*kernel[1]+tmp[8421]*kernel[2]+tmp[8519]*kernel[3]+tmp[8520]*kernel[4]+tmp[8521]*kernel[5]+tmp[8619]*kernel[6]+tmp[8620]*kernel[7]+tmp[8621]*kernel[8];
				ans[8521]<=tmp[8420]*kernel[0]+tmp[8421]*kernel[1]+tmp[8422]*kernel[2]+tmp[8520]*kernel[3]+tmp[8521]*kernel[4]+tmp[8522]*kernel[5]+tmp[8620]*kernel[6]+tmp[8621]*kernel[7]+tmp[8622]*kernel[8];
				ans[8522]<=tmp[8421]*kernel[0]+tmp[8422]*kernel[1]+tmp[8423]*kernel[2]+tmp[8521]*kernel[3]+tmp[8522]*kernel[4]+tmp[8523]*kernel[5]+tmp[8621]*kernel[6]+tmp[8622]*kernel[7]+tmp[8623]*kernel[8];
				ans[8523]<=tmp[8422]*kernel[0]+tmp[8423]*kernel[1]+tmp[8424]*kernel[2]+tmp[8522]*kernel[3]+tmp[8523]*kernel[4]+tmp[8524]*kernel[5]+tmp[8622]*kernel[6]+tmp[8623]*kernel[7]+tmp[8624]*kernel[8];
				ans[8524]<=tmp[8423]*kernel[0]+tmp[8424]*kernel[1]+tmp[8425]*kernel[2]+tmp[8523]*kernel[3]+tmp[8524]*kernel[4]+tmp[8525]*kernel[5]+tmp[8623]*kernel[6]+tmp[8624]*kernel[7]+tmp[8625]*kernel[8];
				ans[8525]<=tmp[8424]*kernel[0]+tmp[8425]*kernel[1]+tmp[8426]*kernel[2]+tmp[8524]*kernel[3]+tmp[8525]*kernel[4]+tmp[8526]*kernel[5]+tmp[8624]*kernel[6]+tmp[8625]*kernel[7]+tmp[8626]*kernel[8];
				ans[8526]<=tmp[8425]*kernel[0]+tmp[8426]*kernel[1]+tmp[8427]*kernel[2]+tmp[8525]*kernel[3]+tmp[8526]*kernel[4]+tmp[8527]*kernel[5]+tmp[8625]*kernel[6]+tmp[8626]*kernel[7]+tmp[8627]*kernel[8];
				ans[8527]<=tmp[8426]*kernel[0]+tmp[8427]*kernel[1]+tmp[8428]*kernel[2]+tmp[8526]*kernel[3]+tmp[8527]*kernel[4]+tmp[8528]*kernel[5]+tmp[8626]*kernel[6]+tmp[8627]*kernel[7]+tmp[8628]*kernel[8];
				ans[8528]<=tmp[8427]*kernel[0]+tmp[8428]*kernel[1]+tmp[8429]*kernel[2]+tmp[8527]*kernel[3]+tmp[8528]*kernel[4]+tmp[8529]*kernel[5]+tmp[8627]*kernel[6]+tmp[8628]*kernel[7]+tmp[8629]*kernel[8];
				ans[8529]<=tmp[8428]*kernel[0]+tmp[8429]*kernel[1]+tmp[8430]*kernel[2]+tmp[8528]*kernel[3]+tmp[8529]*kernel[4]+tmp[8530]*kernel[5]+tmp[8628]*kernel[6]+tmp[8629]*kernel[7]+tmp[8630]*kernel[8];
				ans[8530]<=tmp[8429]*kernel[0]+tmp[8430]*kernel[1]+tmp[8431]*kernel[2]+tmp[8529]*kernel[3]+tmp[8530]*kernel[4]+tmp[8531]*kernel[5]+tmp[8629]*kernel[6]+tmp[8630]*kernel[7]+tmp[8631]*kernel[8];
				ans[8531]<=tmp[8430]*kernel[0]+tmp[8431]*kernel[1]+tmp[8432]*kernel[2]+tmp[8530]*kernel[3]+tmp[8531]*kernel[4]+tmp[8532]*kernel[5]+tmp[8630]*kernel[6]+tmp[8631]*kernel[7]+tmp[8632]*kernel[8];
				ans[8532]<=tmp[8431]*kernel[0]+tmp[8432]*kernel[1]+tmp[8433]*kernel[2]+tmp[8531]*kernel[3]+tmp[8532]*kernel[4]+tmp[8533]*kernel[5]+tmp[8631]*kernel[6]+tmp[8632]*kernel[7]+tmp[8633]*kernel[8];
				ans[8533]<=tmp[8432]*kernel[0]+tmp[8433]*kernel[1]+tmp[8434]*kernel[2]+tmp[8532]*kernel[3]+tmp[8533]*kernel[4]+tmp[8534]*kernel[5]+tmp[8632]*kernel[6]+tmp[8633]*kernel[7]+tmp[8634]*kernel[8];
				ans[8534]<=tmp[8433]*kernel[0]+tmp[8434]*kernel[1]+tmp[8435]*kernel[2]+tmp[8533]*kernel[3]+tmp[8534]*kernel[4]+tmp[8535]*kernel[5]+tmp[8633]*kernel[6]+tmp[8634]*kernel[7]+tmp[8635]*kernel[8];
				ans[8535]<=tmp[8434]*kernel[0]+tmp[8435]*kernel[1]+tmp[8436]*kernel[2]+tmp[8534]*kernel[3]+tmp[8535]*kernel[4]+tmp[8536]*kernel[5]+tmp[8634]*kernel[6]+tmp[8635]*kernel[7]+tmp[8636]*kernel[8];
				ans[8536]<=tmp[8435]*kernel[0]+tmp[8436]*kernel[1]+tmp[8437]*kernel[2]+tmp[8535]*kernel[3]+tmp[8536]*kernel[4]+tmp[8537]*kernel[5]+tmp[8635]*kernel[6]+tmp[8636]*kernel[7]+tmp[8637]*kernel[8];
				ans[8537]<=tmp[8436]*kernel[0]+tmp[8437]*kernel[1]+tmp[8438]*kernel[2]+tmp[8536]*kernel[3]+tmp[8537]*kernel[4]+tmp[8538]*kernel[5]+tmp[8636]*kernel[6]+tmp[8637]*kernel[7]+tmp[8638]*kernel[8];
				ans[8538]<=tmp[8437]*kernel[0]+tmp[8438]*kernel[1]+tmp[8439]*kernel[2]+tmp[8537]*kernel[3]+tmp[8538]*kernel[4]+tmp[8539]*kernel[5]+tmp[8637]*kernel[6]+tmp[8638]*kernel[7]+tmp[8639]*kernel[8];
				ans[8539]<=tmp[8438]*kernel[0]+tmp[8439]*kernel[1]+tmp[8440]*kernel[2]+tmp[8538]*kernel[3]+tmp[8539]*kernel[4]+tmp[8540]*kernel[5]+tmp[8638]*kernel[6]+tmp[8639]*kernel[7]+tmp[8640]*kernel[8];
				ans[8540]<=tmp[8439]*kernel[0]+tmp[8440]*kernel[1]+tmp[8441]*kernel[2]+tmp[8539]*kernel[3]+tmp[8540]*kernel[4]+tmp[8541]*kernel[5]+tmp[8639]*kernel[6]+tmp[8640]*kernel[7]+tmp[8641]*kernel[8];
				ans[8541]<=tmp[8440]*kernel[0]+tmp[8441]*kernel[1]+tmp[8442]*kernel[2]+tmp[8540]*kernel[3]+tmp[8541]*kernel[4]+tmp[8542]*kernel[5]+tmp[8640]*kernel[6]+tmp[8641]*kernel[7]+tmp[8642]*kernel[8];
				ans[8542]<=tmp[8441]*kernel[0]+tmp[8442]*kernel[1]+tmp[8443]*kernel[2]+tmp[8541]*kernel[3]+tmp[8542]*kernel[4]+tmp[8543]*kernel[5]+tmp[8641]*kernel[6]+tmp[8642]*kernel[7]+tmp[8643]*kernel[8];
				ans[8543]<=tmp[8442]*kernel[0]+tmp[8443]*kernel[1]+tmp[8444]*kernel[2]+tmp[8542]*kernel[3]+tmp[8543]*kernel[4]+tmp[8544]*kernel[5]+tmp[8642]*kernel[6]+tmp[8643]*kernel[7]+tmp[8644]*kernel[8];
				ans[8544]<=tmp[8443]*kernel[0]+tmp[8444]*kernel[1]+tmp[8445]*kernel[2]+tmp[8543]*kernel[3]+tmp[8544]*kernel[4]+tmp[8545]*kernel[5]+tmp[8643]*kernel[6]+tmp[8644]*kernel[7]+tmp[8645]*kernel[8];
				ans[8545]<=tmp[8444]*kernel[0]+tmp[8445]*kernel[1]+tmp[8446]*kernel[2]+tmp[8544]*kernel[3]+tmp[8545]*kernel[4]+tmp[8546]*kernel[5]+tmp[8644]*kernel[6]+tmp[8645]*kernel[7]+tmp[8646]*kernel[8];
				ans[8546]<=tmp[8445]*kernel[0]+tmp[8446]*kernel[1]+tmp[8447]*kernel[2]+tmp[8545]*kernel[3]+tmp[8546]*kernel[4]+tmp[8547]*kernel[5]+tmp[8645]*kernel[6]+tmp[8646]*kernel[7]+tmp[8647]*kernel[8];
				ans[8547]<=tmp[8446]*kernel[0]+tmp[8447]*kernel[1]+tmp[8448]*kernel[2]+tmp[8546]*kernel[3]+tmp[8547]*kernel[4]+tmp[8548]*kernel[5]+tmp[8646]*kernel[6]+tmp[8647]*kernel[7]+tmp[8648]*kernel[8];
				ans[8548]<=tmp[8447]*kernel[0]+tmp[8448]*kernel[1]+tmp[8449]*kernel[2]+tmp[8547]*kernel[3]+tmp[8548]*kernel[4]+tmp[8549]*kernel[5]+tmp[8647]*kernel[6]+tmp[8648]*kernel[7]+tmp[8649]*kernel[8];
				ans[8549]<=tmp[8448]*kernel[0]+tmp[8449]*kernel[1]+tmp[8450]*kernel[2]+tmp[8548]*kernel[3]+tmp[8549]*kernel[4]+tmp[8550]*kernel[5]+tmp[8648]*kernel[6]+tmp[8649]*kernel[7]+tmp[8650]*kernel[8];
				ans[8550]<=tmp[8449]*kernel[0]+tmp[8450]*kernel[1]+tmp[8451]*kernel[2]+tmp[8549]*kernel[3]+tmp[8550]*kernel[4]+tmp[8551]*kernel[5]+tmp[8649]*kernel[6]+tmp[8650]*kernel[7]+tmp[8651]*kernel[8];
				ans[8551]<=tmp[8450]*kernel[0]+tmp[8451]*kernel[1]+tmp[8452]*kernel[2]+tmp[8550]*kernel[3]+tmp[8551]*kernel[4]+tmp[8552]*kernel[5]+tmp[8650]*kernel[6]+tmp[8651]*kernel[7]+tmp[8652]*kernel[8];
				ans[8552]<=tmp[8451]*kernel[0]+tmp[8452]*kernel[1]+tmp[8453]*kernel[2]+tmp[8551]*kernel[3]+tmp[8552]*kernel[4]+tmp[8553]*kernel[5]+tmp[8651]*kernel[6]+tmp[8652]*kernel[7]+tmp[8653]*kernel[8];
				ans[8553]<=tmp[8452]*kernel[0]+tmp[8453]*kernel[1]+tmp[8454]*kernel[2]+tmp[8552]*kernel[3]+tmp[8553]*kernel[4]+tmp[8554]*kernel[5]+tmp[8652]*kernel[6]+tmp[8653]*kernel[7]+tmp[8654]*kernel[8];
				ans[8554]<=tmp[8453]*kernel[0]+tmp[8454]*kernel[1]+tmp[8455]*kernel[2]+tmp[8553]*kernel[3]+tmp[8554]*kernel[4]+tmp[8555]*kernel[5]+tmp[8653]*kernel[6]+tmp[8654]*kernel[7]+tmp[8655]*kernel[8];
				ans[8555]<=tmp[8454]*kernel[0]+tmp[8455]*kernel[1]+tmp[8456]*kernel[2]+tmp[8554]*kernel[3]+tmp[8555]*kernel[4]+tmp[8556]*kernel[5]+tmp[8654]*kernel[6]+tmp[8655]*kernel[7]+tmp[8656]*kernel[8];
				ans[8556]<=tmp[8455]*kernel[0]+tmp[8456]*kernel[1]+tmp[8457]*kernel[2]+tmp[8555]*kernel[3]+tmp[8556]*kernel[4]+tmp[8557]*kernel[5]+tmp[8655]*kernel[6]+tmp[8656]*kernel[7]+tmp[8657]*kernel[8];
				ans[8557]<=tmp[8456]*kernel[0]+tmp[8457]*kernel[1]+tmp[8458]*kernel[2]+tmp[8556]*kernel[3]+tmp[8557]*kernel[4]+tmp[8558]*kernel[5]+tmp[8656]*kernel[6]+tmp[8657]*kernel[7]+tmp[8658]*kernel[8];
				ans[8558]<=tmp[8457]*kernel[0]+tmp[8458]*kernel[1]+tmp[8459]*kernel[2]+tmp[8557]*kernel[3]+tmp[8558]*kernel[4]+tmp[8559]*kernel[5]+tmp[8657]*kernel[6]+tmp[8658]*kernel[7]+tmp[8659]*kernel[8];
				ans[8559]<=tmp[8458]*kernel[0]+tmp[8459]*kernel[1]+tmp[8460]*kernel[2]+tmp[8558]*kernel[3]+tmp[8559]*kernel[4]+tmp[8560]*kernel[5]+tmp[8658]*kernel[6]+tmp[8659]*kernel[7]+tmp[8660]*kernel[8];
				ans[8560]<=tmp[8459]*kernel[0]+tmp[8460]*kernel[1]+tmp[8461]*kernel[2]+tmp[8559]*kernel[3]+tmp[8560]*kernel[4]+tmp[8561]*kernel[5]+tmp[8659]*kernel[6]+tmp[8660]*kernel[7]+tmp[8661]*kernel[8];
				ans[8561]<=tmp[8460]*kernel[0]+tmp[8461]*kernel[1]+tmp[8462]*kernel[2]+tmp[8560]*kernel[3]+tmp[8561]*kernel[4]+tmp[8562]*kernel[5]+tmp[8660]*kernel[6]+tmp[8661]*kernel[7]+tmp[8662]*kernel[8];
				ans[8562]<=tmp[8461]*kernel[0]+tmp[8462]*kernel[1]+tmp[8463]*kernel[2]+tmp[8561]*kernel[3]+tmp[8562]*kernel[4]+tmp[8563]*kernel[5]+tmp[8661]*kernel[6]+tmp[8662]*kernel[7]+tmp[8663]*kernel[8];
				ans[8563]<=tmp[8462]*kernel[0]+tmp[8463]*kernel[1]+tmp[8464]*kernel[2]+tmp[8562]*kernel[3]+tmp[8563]*kernel[4]+tmp[8564]*kernel[5]+tmp[8662]*kernel[6]+tmp[8663]*kernel[7]+tmp[8664]*kernel[8];
				ans[8564]<=tmp[8463]*kernel[0]+tmp[8464]*kernel[1]+tmp[8465]*kernel[2]+tmp[8563]*kernel[3]+tmp[8564]*kernel[4]+tmp[8565]*kernel[5]+tmp[8663]*kernel[6]+tmp[8664]*kernel[7]+tmp[8665]*kernel[8];
				ans[8565]<=tmp[8464]*kernel[0]+tmp[8465]*kernel[1]+tmp[8466]*kernel[2]+tmp[8564]*kernel[3]+tmp[8565]*kernel[4]+tmp[8566]*kernel[5]+tmp[8664]*kernel[6]+tmp[8665]*kernel[7]+tmp[8666]*kernel[8];
				ans[8566]<=tmp[8465]*kernel[0]+tmp[8466]*kernel[1]+tmp[8467]*kernel[2]+tmp[8565]*kernel[3]+tmp[8566]*kernel[4]+tmp[8567]*kernel[5]+tmp[8665]*kernel[6]+tmp[8666]*kernel[7]+tmp[8667]*kernel[8];
				ans[8567]<=tmp[8466]*kernel[0]+tmp[8467]*kernel[1]+tmp[8468]*kernel[2]+tmp[8566]*kernel[3]+tmp[8567]*kernel[4]+tmp[8568]*kernel[5]+tmp[8666]*kernel[6]+tmp[8667]*kernel[7]+tmp[8668]*kernel[8];
				ans[8568]<=tmp[8467]*kernel[0]+tmp[8468]*kernel[1]+tmp[8469]*kernel[2]+tmp[8567]*kernel[3]+tmp[8568]*kernel[4]+tmp[8569]*kernel[5]+tmp[8667]*kernel[6]+tmp[8668]*kernel[7]+tmp[8669]*kernel[8];
				ans[8569]<=tmp[8468]*kernel[0]+tmp[8469]*kernel[1]+tmp[8470]*kernel[2]+tmp[8568]*kernel[3]+tmp[8569]*kernel[4]+tmp[8570]*kernel[5]+tmp[8668]*kernel[6]+tmp[8669]*kernel[7]+tmp[8670]*kernel[8];
				ans[8570]<=tmp[8469]*kernel[0]+tmp[8470]*kernel[1]+tmp[8471]*kernel[2]+tmp[8569]*kernel[3]+tmp[8570]*kernel[4]+tmp[8571]*kernel[5]+tmp[8669]*kernel[6]+tmp[8670]*kernel[7]+tmp[8671]*kernel[8];
				ans[8571]<=tmp[8470]*kernel[0]+tmp[8471]*kernel[1]+tmp[8472]*kernel[2]+tmp[8570]*kernel[3]+tmp[8571]*kernel[4]+tmp[8572]*kernel[5]+tmp[8670]*kernel[6]+tmp[8671]*kernel[7]+tmp[8672]*kernel[8];
				ans[8572]<=tmp[8471]*kernel[0]+tmp[8472]*kernel[1]+tmp[8473]*kernel[2]+tmp[8571]*kernel[3]+tmp[8572]*kernel[4]+tmp[8573]*kernel[5]+tmp[8671]*kernel[6]+tmp[8672]*kernel[7]+tmp[8673]*kernel[8];
				ans[8573]<=tmp[8472]*kernel[0]+tmp[8473]*kernel[1]+tmp[8474]*kernel[2]+tmp[8572]*kernel[3]+tmp[8573]*kernel[4]+tmp[8574]*kernel[5]+tmp[8672]*kernel[6]+tmp[8673]*kernel[7]+tmp[8674]*kernel[8];
				ans[8574]<=tmp[8473]*kernel[0]+tmp[8474]*kernel[1]+tmp[8475]*kernel[2]+tmp[8573]*kernel[3]+tmp[8574]*kernel[4]+tmp[8575]*kernel[5]+tmp[8673]*kernel[6]+tmp[8674]*kernel[7]+tmp[8675]*kernel[8];
				ans[8575]<=tmp[8474]*kernel[0]+tmp[8475]*kernel[1]+tmp[8476]*kernel[2]+tmp[8574]*kernel[3]+tmp[8575]*kernel[4]+tmp[8576]*kernel[5]+tmp[8674]*kernel[6]+tmp[8675]*kernel[7]+tmp[8676]*kernel[8];
				ans[8576]<=tmp[8475]*kernel[0]+tmp[8476]*kernel[1]+tmp[8477]*kernel[2]+tmp[8575]*kernel[3]+tmp[8576]*kernel[4]+tmp[8577]*kernel[5]+tmp[8675]*kernel[6]+tmp[8676]*kernel[7]+tmp[8677]*kernel[8];
				ans[8577]<=tmp[8476]*kernel[0]+tmp[8477]*kernel[1]+tmp[8478]*kernel[2]+tmp[8576]*kernel[3]+tmp[8577]*kernel[4]+tmp[8578]*kernel[5]+tmp[8676]*kernel[6]+tmp[8677]*kernel[7]+tmp[8678]*kernel[8];
				ans[8578]<=tmp[8477]*kernel[0]+tmp[8478]*kernel[1]+tmp[8479]*kernel[2]+tmp[8577]*kernel[3]+tmp[8578]*kernel[4]+tmp[8579]*kernel[5]+tmp[8677]*kernel[6]+tmp[8678]*kernel[7]+tmp[8679]*kernel[8];
				ans[8579]<=tmp[8478]*kernel[0]+tmp[8479]*kernel[1]+tmp[8480]*kernel[2]+tmp[8578]*kernel[3]+tmp[8579]*kernel[4]+tmp[8580]*kernel[5]+tmp[8678]*kernel[6]+tmp[8679]*kernel[7]+tmp[8680]*kernel[8];
				ans[8580]<=tmp[8479]*kernel[0]+tmp[8480]*kernel[1]+tmp[8481]*kernel[2]+tmp[8579]*kernel[3]+tmp[8580]*kernel[4]+tmp[8581]*kernel[5]+tmp[8679]*kernel[6]+tmp[8680]*kernel[7]+tmp[8681]*kernel[8];
				ans[8581]<=tmp[8480]*kernel[0]+tmp[8481]*kernel[1]+tmp[8482]*kernel[2]+tmp[8580]*kernel[3]+tmp[8581]*kernel[4]+tmp[8582]*kernel[5]+tmp[8680]*kernel[6]+tmp[8681]*kernel[7]+tmp[8682]*kernel[8];
				ans[8582]<=tmp[8481]*kernel[0]+tmp[8482]*kernel[1]+tmp[8483]*kernel[2]+tmp[8581]*kernel[3]+tmp[8582]*kernel[4]+tmp[8583]*kernel[5]+tmp[8681]*kernel[6]+tmp[8682]*kernel[7]+tmp[8683]*kernel[8];
				ans[8583]<=tmp[8482]*kernel[0]+tmp[8483]*kernel[1]+tmp[8484]*kernel[2]+tmp[8582]*kernel[3]+tmp[8583]*kernel[4]+tmp[8584]*kernel[5]+tmp[8682]*kernel[6]+tmp[8683]*kernel[7]+tmp[8684]*kernel[8];
				ans[8584]<=tmp[8483]*kernel[0]+tmp[8484]*kernel[1]+tmp[8485]*kernel[2]+tmp[8583]*kernel[3]+tmp[8584]*kernel[4]+tmp[8585]*kernel[5]+tmp[8683]*kernel[6]+tmp[8684]*kernel[7]+tmp[8685]*kernel[8];
				ans[8585]<=tmp[8484]*kernel[0]+tmp[8485]*kernel[1]+tmp[8486]*kernel[2]+tmp[8584]*kernel[3]+tmp[8585]*kernel[4]+tmp[8586]*kernel[5]+tmp[8684]*kernel[6]+tmp[8685]*kernel[7]+tmp[8686]*kernel[8];
				ans[8586]<=tmp[8485]*kernel[0]+tmp[8486]*kernel[1]+tmp[8487]*kernel[2]+tmp[8585]*kernel[3]+tmp[8586]*kernel[4]+tmp[8587]*kernel[5]+tmp[8685]*kernel[6]+tmp[8686]*kernel[7]+tmp[8687]*kernel[8];
				ans[8587]<=tmp[8486]*kernel[0]+tmp[8487]*kernel[1]+tmp[8488]*kernel[2]+tmp[8586]*kernel[3]+tmp[8587]*kernel[4]+tmp[8588]*kernel[5]+tmp[8686]*kernel[6]+tmp[8687]*kernel[7]+tmp[8688]*kernel[8];
				ans[8588]<=tmp[8487]*kernel[0]+tmp[8488]*kernel[1]+tmp[8489]*kernel[2]+tmp[8587]*kernel[3]+tmp[8588]*kernel[4]+tmp[8589]*kernel[5]+tmp[8687]*kernel[6]+tmp[8688]*kernel[7]+tmp[8689]*kernel[8];
				ans[8589]<=tmp[8488]*kernel[0]+tmp[8489]*kernel[1]+tmp[8490]*kernel[2]+tmp[8588]*kernel[3]+tmp[8589]*kernel[4]+tmp[8590]*kernel[5]+tmp[8688]*kernel[6]+tmp[8689]*kernel[7]+tmp[8690]*kernel[8];
				ans[8590]<=tmp[8489]*kernel[0]+tmp[8490]*kernel[1]+tmp[8491]*kernel[2]+tmp[8589]*kernel[3]+tmp[8590]*kernel[4]+tmp[8591]*kernel[5]+tmp[8689]*kernel[6]+tmp[8690]*kernel[7]+tmp[8691]*kernel[8];
				ans[8591]<=tmp[8490]*kernel[0]+tmp[8491]*kernel[1]+tmp[8492]*kernel[2]+tmp[8590]*kernel[3]+tmp[8591]*kernel[4]+tmp[8592]*kernel[5]+tmp[8690]*kernel[6]+tmp[8691]*kernel[7]+tmp[8692]*kernel[8];
				ans[8592]<=tmp[8491]*kernel[0]+tmp[8492]*kernel[1]+tmp[8493]*kernel[2]+tmp[8591]*kernel[3]+tmp[8592]*kernel[4]+tmp[8593]*kernel[5]+tmp[8691]*kernel[6]+tmp[8692]*kernel[7]+tmp[8693]*kernel[8];
				ans[8593]<=tmp[8492]*kernel[0]+tmp[8493]*kernel[1]+tmp[8494]*kernel[2]+tmp[8592]*kernel[3]+tmp[8593]*kernel[4]+tmp[8594]*kernel[5]+tmp[8692]*kernel[6]+tmp[8693]*kernel[7]+tmp[8694]*kernel[8];
				ans[8594]<=tmp[8493]*kernel[0]+tmp[8494]*kernel[1]+tmp[8495]*kernel[2]+tmp[8593]*kernel[3]+tmp[8594]*kernel[4]+tmp[8595]*kernel[5]+tmp[8693]*kernel[6]+tmp[8694]*kernel[7]+tmp[8695]*kernel[8];
				ans[8595]<=tmp[8494]*kernel[0]+tmp[8495]*kernel[1]+tmp[8496]*kernel[2]+tmp[8594]*kernel[3]+tmp[8595]*kernel[4]+tmp[8596]*kernel[5]+tmp[8694]*kernel[6]+tmp[8695]*kernel[7]+tmp[8696]*kernel[8];
				ans[8596]<=tmp[8495]*kernel[0]+tmp[8496]*kernel[1]+tmp[8497]*kernel[2]+tmp[8595]*kernel[3]+tmp[8596]*kernel[4]+tmp[8597]*kernel[5]+tmp[8695]*kernel[6]+tmp[8696]*kernel[7]+tmp[8697]*kernel[8];
				ans[8597]<=tmp[8496]*kernel[0]+tmp[8497]*kernel[1]+tmp[8498]*kernel[2]+tmp[8596]*kernel[3]+tmp[8597]*kernel[4]+tmp[8598]*kernel[5]+tmp[8696]*kernel[6]+tmp[8697]*kernel[7]+tmp[8698]*kernel[8];
				ans[8598]<=tmp[8497]*kernel[0]+tmp[8498]*kernel[1]+tmp[8499]*kernel[2]+tmp[8597]*kernel[3]+tmp[8598]*kernel[4]+tmp[8599]*kernel[5]+tmp[8697]*kernel[6]+tmp[8698]*kernel[7]+tmp[8699]*kernel[8];
				ans[8599]<=tmp[8498]*kernel[0]+tmp[8499]*kernel[1]+tmp[8598]*kernel[3]+tmp[8599]*kernel[4]+tmp[8698]*kernel[6]+tmp[8699]*kernel[7];
				ans[8600]<=tmp[8500]*kernel[1]+tmp[8501]*kernel[2]+tmp[8600]*kernel[4]+tmp[8601]*kernel[5]+tmp[8700]*kernel[7]+tmp[8701]*kernel[8];
				ans[8601]<=tmp[8500]*kernel[0]+tmp[8501]*kernel[1]+tmp[8502]*kernel[2]+tmp[8600]*kernel[3]+tmp[8601]*kernel[4]+tmp[8602]*kernel[5]+tmp[8700]*kernel[6]+tmp[8701]*kernel[7]+tmp[8702]*kernel[8];
				ans[8602]<=tmp[8501]*kernel[0]+tmp[8502]*kernel[1]+tmp[8503]*kernel[2]+tmp[8601]*kernel[3]+tmp[8602]*kernel[4]+tmp[8603]*kernel[5]+tmp[8701]*kernel[6]+tmp[8702]*kernel[7]+tmp[8703]*kernel[8];
				ans[8603]<=tmp[8502]*kernel[0]+tmp[8503]*kernel[1]+tmp[8504]*kernel[2]+tmp[8602]*kernel[3]+tmp[8603]*kernel[4]+tmp[8604]*kernel[5]+tmp[8702]*kernel[6]+tmp[8703]*kernel[7]+tmp[8704]*kernel[8];
				ans[8604]<=tmp[8503]*kernel[0]+tmp[8504]*kernel[1]+tmp[8505]*kernel[2]+tmp[8603]*kernel[3]+tmp[8604]*kernel[4]+tmp[8605]*kernel[5]+tmp[8703]*kernel[6]+tmp[8704]*kernel[7]+tmp[8705]*kernel[8];
				ans[8605]<=tmp[8504]*kernel[0]+tmp[8505]*kernel[1]+tmp[8506]*kernel[2]+tmp[8604]*kernel[3]+tmp[8605]*kernel[4]+tmp[8606]*kernel[5]+tmp[8704]*kernel[6]+tmp[8705]*kernel[7]+tmp[8706]*kernel[8];
				ans[8606]<=tmp[8505]*kernel[0]+tmp[8506]*kernel[1]+tmp[8507]*kernel[2]+tmp[8605]*kernel[3]+tmp[8606]*kernel[4]+tmp[8607]*kernel[5]+tmp[8705]*kernel[6]+tmp[8706]*kernel[7]+tmp[8707]*kernel[8];
				ans[8607]<=tmp[8506]*kernel[0]+tmp[8507]*kernel[1]+tmp[8508]*kernel[2]+tmp[8606]*kernel[3]+tmp[8607]*kernel[4]+tmp[8608]*kernel[5]+tmp[8706]*kernel[6]+tmp[8707]*kernel[7]+tmp[8708]*kernel[8];
				ans[8608]<=tmp[8507]*kernel[0]+tmp[8508]*kernel[1]+tmp[8509]*kernel[2]+tmp[8607]*kernel[3]+tmp[8608]*kernel[4]+tmp[8609]*kernel[5]+tmp[8707]*kernel[6]+tmp[8708]*kernel[7]+tmp[8709]*kernel[8];
				ans[8609]<=tmp[8508]*kernel[0]+tmp[8509]*kernel[1]+tmp[8510]*kernel[2]+tmp[8608]*kernel[3]+tmp[8609]*kernel[4]+tmp[8610]*kernel[5]+tmp[8708]*kernel[6]+tmp[8709]*kernel[7]+tmp[8710]*kernel[8];
				ans[8610]<=tmp[8509]*kernel[0]+tmp[8510]*kernel[1]+tmp[8511]*kernel[2]+tmp[8609]*kernel[3]+tmp[8610]*kernel[4]+tmp[8611]*kernel[5]+tmp[8709]*kernel[6]+tmp[8710]*kernel[7]+tmp[8711]*kernel[8];
				ans[8611]<=tmp[8510]*kernel[0]+tmp[8511]*kernel[1]+tmp[8512]*kernel[2]+tmp[8610]*kernel[3]+tmp[8611]*kernel[4]+tmp[8612]*kernel[5]+tmp[8710]*kernel[6]+tmp[8711]*kernel[7]+tmp[8712]*kernel[8];
				ans[8612]<=tmp[8511]*kernel[0]+tmp[8512]*kernel[1]+tmp[8513]*kernel[2]+tmp[8611]*kernel[3]+tmp[8612]*kernel[4]+tmp[8613]*kernel[5]+tmp[8711]*kernel[6]+tmp[8712]*kernel[7]+tmp[8713]*kernel[8];
				ans[8613]<=tmp[8512]*kernel[0]+tmp[8513]*kernel[1]+tmp[8514]*kernel[2]+tmp[8612]*kernel[3]+tmp[8613]*kernel[4]+tmp[8614]*kernel[5]+tmp[8712]*kernel[6]+tmp[8713]*kernel[7]+tmp[8714]*kernel[8];
				ans[8614]<=tmp[8513]*kernel[0]+tmp[8514]*kernel[1]+tmp[8515]*kernel[2]+tmp[8613]*kernel[3]+tmp[8614]*kernel[4]+tmp[8615]*kernel[5]+tmp[8713]*kernel[6]+tmp[8714]*kernel[7]+tmp[8715]*kernel[8];
				ans[8615]<=tmp[8514]*kernel[0]+tmp[8515]*kernel[1]+tmp[8516]*kernel[2]+tmp[8614]*kernel[3]+tmp[8615]*kernel[4]+tmp[8616]*kernel[5]+tmp[8714]*kernel[6]+tmp[8715]*kernel[7]+tmp[8716]*kernel[8];
				ans[8616]<=tmp[8515]*kernel[0]+tmp[8516]*kernel[1]+tmp[8517]*kernel[2]+tmp[8615]*kernel[3]+tmp[8616]*kernel[4]+tmp[8617]*kernel[5]+tmp[8715]*kernel[6]+tmp[8716]*kernel[7]+tmp[8717]*kernel[8];
				ans[8617]<=tmp[8516]*kernel[0]+tmp[8517]*kernel[1]+tmp[8518]*kernel[2]+tmp[8616]*kernel[3]+tmp[8617]*kernel[4]+tmp[8618]*kernel[5]+tmp[8716]*kernel[6]+tmp[8717]*kernel[7]+tmp[8718]*kernel[8];
				ans[8618]<=tmp[8517]*kernel[0]+tmp[8518]*kernel[1]+tmp[8519]*kernel[2]+tmp[8617]*kernel[3]+tmp[8618]*kernel[4]+tmp[8619]*kernel[5]+tmp[8717]*kernel[6]+tmp[8718]*kernel[7]+tmp[8719]*kernel[8];
				ans[8619]<=tmp[8518]*kernel[0]+tmp[8519]*kernel[1]+tmp[8520]*kernel[2]+tmp[8618]*kernel[3]+tmp[8619]*kernel[4]+tmp[8620]*kernel[5]+tmp[8718]*kernel[6]+tmp[8719]*kernel[7]+tmp[8720]*kernel[8];
				ans[8620]<=tmp[8519]*kernel[0]+tmp[8520]*kernel[1]+tmp[8521]*kernel[2]+tmp[8619]*kernel[3]+tmp[8620]*kernel[4]+tmp[8621]*kernel[5]+tmp[8719]*kernel[6]+tmp[8720]*kernel[7]+tmp[8721]*kernel[8];
				ans[8621]<=tmp[8520]*kernel[0]+tmp[8521]*kernel[1]+tmp[8522]*kernel[2]+tmp[8620]*kernel[3]+tmp[8621]*kernel[4]+tmp[8622]*kernel[5]+tmp[8720]*kernel[6]+tmp[8721]*kernel[7]+tmp[8722]*kernel[8];
				ans[8622]<=tmp[8521]*kernel[0]+tmp[8522]*kernel[1]+tmp[8523]*kernel[2]+tmp[8621]*kernel[3]+tmp[8622]*kernel[4]+tmp[8623]*kernel[5]+tmp[8721]*kernel[6]+tmp[8722]*kernel[7]+tmp[8723]*kernel[8];
				ans[8623]<=tmp[8522]*kernel[0]+tmp[8523]*kernel[1]+tmp[8524]*kernel[2]+tmp[8622]*kernel[3]+tmp[8623]*kernel[4]+tmp[8624]*kernel[5]+tmp[8722]*kernel[6]+tmp[8723]*kernel[7]+tmp[8724]*kernel[8];
				ans[8624]<=tmp[8523]*kernel[0]+tmp[8524]*kernel[1]+tmp[8525]*kernel[2]+tmp[8623]*kernel[3]+tmp[8624]*kernel[4]+tmp[8625]*kernel[5]+tmp[8723]*kernel[6]+tmp[8724]*kernel[7]+tmp[8725]*kernel[8];
				ans[8625]<=tmp[8524]*kernel[0]+tmp[8525]*kernel[1]+tmp[8526]*kernel[2]+tmp[8624]*kernel[3]+tmp[8625]*kernel[4]+tmp[8626]*kernel[5]+tmp[8724]*kernel[6]+tmp[8725]*kernel[7]+tmp[8726]*kernel[8];
				ans[8626]<=tmp[8525]*kernel[0]+tmp[8526]*kernel[1]+tmp[8527]*kernel[2]+tmp[8625]*kernel[3]+tmp[8626]*kernel[4]+tmp[8627]*kernel[5]+tmp[8725]*kernel[6]+tmp[8726]*kernel[7]+tmp[8727]*kernel[8];
				ans[8627]<=tmp[8526]*kernel[0]+tmp[8527]*kernel[1]+tmp[8528]*kernel[2]+tmp[8626]*kernel[3]+tmp[8627]*kernel[4]+tmp[8628]*kernel[5]+tmp[8726]*kernel[6]+tmp[8727]*kernel[7]+tmp[8728]*kernel[8];
				ans[8628]<=tmp[8527]*kernel[0]+tmp[8528]*kernel[1]+tmp[8529]*kernel[2]+tmp[8627]*kernel[3]+tmp[8628]*kernel[4]+tmp[8629]*kernel[5]+tmp[8727]*kernel[6]+tmp[8728]*kernel[7]+tmp[8729]*kernel[8];
				ans[8629]<=tmp[8528]*kernel[0]+tmp[8529]*kernel[1]+tmp[8530]*kernel[2]+tmp[8628]*kernel[3]+tmp[8629]*kernel[4]+tmp[8630]*kernel[5]+tmp[8728]*kernel[6]+tmp[8729]*kernel[7]+tmp[8730]*kernel[8];
				ans[8630]<=tmp[8529]*kernel[0]+tmp[8530]*kernel[1]+tmp[8531]*kernel[2]+tmp[8629]*kernel[3]+tmp[8630]*kernel[4]+tmp[8631]*kernel[5]+tmp[8729]*kernel[6]+tmp[8730]*kernel[7]+tmp[8731]*kernel[8];
				ans[8631]<=tmp[8530]*kernel[0]+tmp[8531]*kernel[1]+tmp[8532]*kernel[2]+tmp[8630]*kernel[3]+tmp[8631]*kernel[4]+tmp[8632]*kernel[5]+tmp[8730]*kernel[6]+tmp[8731]*kernel[7]+tmp[8732]*kernel[8];
				ans[8632]<=tmp[8531]*kernel[0]+tmp[8532]*kernel[1]+tmp[8533]*kernel[2]+tmp[8631]*kernel[3]+tmp[8632]*kernel[4]+tmp[8633]*kernel[5]+tmp[8731]*kernel[6]+tmp[8732]*kernel[7]+tmp[8733]*kernel[8];
				ans[8633]<=tmp[8532]*kernel[0]+tmp[8533]*kernel[1]+tmp[8534]*kernel[2]+tmp[8632]*kernel[3]+tmp[8633]*kernel[4]+tmp[8634]*kernel[5]+tmp[8732]*kernel[6]+tmp[8733]*kernel[7]+tmp[8734]*kernel[8];
				ans[8634]<=tmp[8533]*kernel[0]+tmp[8534]*kernel[1]+tmp[8535]*kernel[2]+tmp[8633]*kernel[3]+tmp[8634]*kernel[4]+tmp[8635]*kernel[5]+tmp[8733]*kernel[6]+tmp[8734]*kernel[7]+tmp[8735]*kernel[8];
				ans[8635]<=tmp[8534]*kernel[0]+tmp[8535]*kernel[1]+tmp[8536]*kernel[2]+tmp[8634]*kernel[3]+tmp[8635]*kernel[4]+tmp[8636]*kernel[5]+tmp[8734]*kernel[6]+tmp[8735]*kernel[7]+tmp[8736]*kernel[8];
				ans[8636]<=tmp[8535]*kernel[0]+tmp[8536]*kernel[1]+tmp[8537]*kernel[2]+tmp[8635]*kernel[3]+tmp[8636]*kernel[4]+tmp[8637]*kernel[5]+tmp[8735]*kernel[6]+tmp[8736]*kernel[7]+tmp[8737]*kernel[8];
				ans[8637]<=tmp[8536]*kernel[0]+tmp[8537]*kernel[1]+tmp[8538]*kernel[2]+tmp[8636]*kernel[3]+tmp[8637]*kernel[4]+tmp[8638]*kernel[5]+tmp[8736]*kernel[6]+tmp[8737]*kernel[7]+tmp[8738]*kernel[8];
				ans[8638]<=tmp[8537]*kernel[0]+tmp[8538]*kernel[1]+tmp[8539]*kernel[2]+tmp[8637]*kernel[3]+tmp[8638]*kernel[4]+tmp[8639]*kernel[5]+tmp[8737]*kernel[6]+tmp[8738]*kernel[7]+tmp[8739]*kernel[8];
				ans[8639]<=tmp[8538]*kernel[0]+tmp[8539]*kernel[1]+tmp[8540]*kernel[2]+tmp[8638]*kernel[3]+tmp[8639]*kernel[4]+tmp[8640]*kernel[5]+tmp[8738]*kernel[6]+tmp[8739]*kernel[7]+tmp[8740]*kernel[8];
				ans[8640]<=tmp[8539]*kernel[0]+tmp[8540]*kernel[1]+tmp[8541]*kernel[2]+tmp[8639]*kernel[3]+tmp[8640]*kernel[4]+tmp[8641]*kernel[5]+tmp[8739]*kernel[6]+tmp[8740]*kernel[7]+tmp[8741]*kernel[8];
				ans[8641]<=tmp[8540]*kernel[0]+tmp[8541]*kernel[1]+tmp[8542]*kernel[2]+tmp[8640]*kernel[3]+tmp[8641]*kernel[4]+tmp[8642]*kernel[5]+tmp[8740]*kernel[6]+tmp[8741]*kernel[7]+tmp[8742]*kernel[8];
				ans[8642]<=tmp[8541]*kernel[0]+tmp[8542]*kernel[1]+tmp[8543]*kernel[2]+tmp[8641]*kernel[3]+tmp[8642]*kernel[4]+tmp[8643]*kernel[5]+tmp[8741]*kernel[6]+tmp[8742]*kernel[7]+tmp[8743]*kernel[8];
				ans[8643]<=tmp[8542]*kernel[0]+tmp[8543]*kernel[1]+tmp[8544]*kernel[2]+tmp[8642]*kernel[3]+tmp[8643]*kernel[4]+tmp[8644]*kernel[5]+tmp[8742]*kernel[6]+tmp[8743]*kernel[7]+tmp[8744]*kernel[8];
				ans[8644]<=tmp[8543]*kernel[0]+tmp[8544]*kernel[1]+tmp[8545]*kernel[2]+tmp[8643]*kernel[3]+tmp[8644]*kernel[4]+tmp[8645]*kernel[5]+tmp[8743]*kernel[6]+tmp[8744]*kernel[7]+tmp[8745]*kernel[8];
				ans[8645]<=tmp[8544]*kernel[0]+tmp[8545]*kernel[1]+tmp[8546]*kernel[2]+tmp[8644]*kernel[3]+tmp[8645]*kernel[4]+tmp[8646]*kernel[5]+tmp[8744]*kernel[6]+tmp[8745]*kernel[7]+tmp[8746]*kernel[8];
				ans[8646]<=tmp[8545]*kernel[0]+tmp[8546]*kernel[1]+tmp[8547]*kernel[2]+tmp[8645]*kernel[3]+tmp[8646]*kernel[4]+tmp[8647]*kernel[5]+tmp[8745]*kernel[6]+tmp[8746]*kernel[7]+tmp[8747]*kernel[8];
				ans[8647]<=tmp[8546]*kernel[0]+tmp[8547]*kernel[1]+tmp[8548]*kernel[2]+tmp[8646]*kernel[3]+tmp[8647]*kernel[4]+tmp[8648]*kernel[5]+tmp[8746]*kernel[6]+tmp[8747]*kernel[7]+tmp[8748]*kernel[8];
				ans[8648]<=tmp[8547]*kernel[0]+tmp[8548]*kernel[1]+tmp[8549]*kernel[2]+tmp[8647]*kernel[3]+tmp[8648]*kernel[4]+tmp[8649]*kernel[5]+tmp[8747]*kernel[6]+tmp[8748]*kernel[7]+tmp[8749]*kernel[8];
				ans[8649]<=tmp[8548]*kernel[0]+tmp[8549]*kernel[1]+tmp[8550]*kernel[2]+tmp[8648]*kernel[3]+tmp[8649]*kernel[4]+tmp[8650]*kernel[5]+tmp[8748]*kernel[6]+tmp[8749]*kernel[7]+tmp[8750]*kernel[8];
				ans[8650]<=tmp[8549]*kernel[0]+tmp[8550]*kernel[1]+tmp[8551]*kernel[2]+tmp[8649]*kernel[3]+tmp[8650]*kernel[4]+tmp[8651]*kernel[5]+tmp[8749]*kernel[6]+tmp[8750]*kernel[7]+tmp[8751]*kernel[8];
				ans[8651]<=tmp[8550]*kernel[0]+tmp[8551]*kernel[1]+tmp[8552]*kernel[2]+tmp[8650]*kernel[3]+tmp[8651]*kernel[4]+tmp[8652]*kernel[5]+tmp[8750]*kernel[6]+tmp[8751]*kernel[7]+tmp[8752]*kernel[8];
				ans[8652]<=tmp[8551]*kernel[0]+tmp[8552]*kernel[1]+tmp[8553]*kernel[2]+tmp[8651]*kernel[3]+tmp[8652]*kernel[4]+tmp[8653]*kernel[5]+tmp[8751]*kernel[6]+tmp[8752]*kernel[7]+tmp[8753]*kernel[8];
				ans[8653]<=tmp[8552]*kernel[0]+tmp[8553]*kernel[1]+tmp[8554]*kernel[2]+tmp[8652]*kernel[3]+tmp[8653]*kernel[4]+tmp[8654]*kernel[5]+tmp[8752]*kernel[6]+tmp[8753]*kernel[7]+tmp[8754]*kernel[8];
				ans[8654]<=tmp[8553]*kernel[0]+tmp[8554]*kernel[1]+tmp[8555]*kernel[2]+tmp[8653]*kernel[3]+tmp[8654]*kernel[4]+tmp[8655]*kernel[5]+tmp[8753]*kernel[6]+tmp[8754]*kernel[7]+tmp[8755]*kernel[8];
				ans[8655]<=tmp[8554]*kernel[0]+tmp[8555]*kernel[1]+tmp[8556]*kernel[2]+tmp[8654]*kernel[3]+tmp[8655]*kernel[4]+tmp[8656]*kernel[5]+tmp[8754]*kernel[6]+tmp[8755]*kernel[7]+tmp[8756]*kernel[8];
				ans[8656]<=tmp[8555]*kernel[0]+tmp[8556]*kernel[1]+tmp[8557]*kernel[2]+tmp[8655]*kernel[3]+tmp[8656]*kernel[4]+tmp[8657]*kernel[5]+tmp[8755]*kernel[6]+tmp[8756]*kernel[7]+tmp[8757]*kernel[8];
				ans[8657]<=tmp[8556]*kernel[0]+tmp[8557]*kernel[1]+tmp[8558]*kernel[2]+tmp[8656]*kernel[3]+tmp[8657]*kernel[4]+tmp[8658]*kernel[5]+tmp[8756]*kernel[6]+tmp[8757]*kernel[7]+tmp[8758]*kernel[8];
				ans[8658]<=tmp[8557]*kernel[0]+tmp[8558]*kernel[1]+tmp[8559]*kernel[2]+tmp[8657]*kernel[3]+tmp[8658]*kernel[4]+tmp[8659]*kernel[5]+tmp[8757]*kernel[6]+tmp[8758]*kernel[7]+tmp[8759]*kernel[8];
				ans[8659]<=tmp[8558]*kernel[0]+tmp[8559]*kernel[1]+tmp[8560]*kernel[2]+tmp[8658]*kernel[3]+tmp[8659]*kernel[4]+tmp[8660]*kernel[5]+tmp[8758]*kernel[6]+tmp[8759]*kernel[7]+tmp[8760]*kernel[8];
				ans[8660]<=tmp[8559]*kernel[0]+tmp[8560]*kernel[1]+tmp[8561]*kernel[2]+tmp[8659]*kernel[3]+tmp[8660]*kernel[4]+tmp[8661]*kernel[5]+tmp[8759]*kernel[6]+tmp[8760]*kernel[7]+tmp[8761]*kernel[8];
				ans[8661]<=tmp[8560]*kernel[0]+tmp[8561]*kernel[1]+tmp[8562]*kernel[2]+tmp[8660]*kernel[3]+tmp[8661]*kernel[4]+tmp[8662]*kernel[5]+tmp[8760]*kernel[6]+tmp[8761]*kernel[7]+tmp[8762]*kernel[8];
				ans[8662]<=tmp[8561]*kernel[0]+tmp[8562]*kernel[1]+tmp[8563]*kernel[2]+tmp[8661]*kernel[3]+tmp[8662]*kernel[4]+tmp[8663]*kernel[5]+tmp[8761]*kernel[6]+tmp[8762]*kernel[7]+tmp[8763]*kernel[8];
				ans[8663]<=tmp[8562]*kernel[0]+tmp[8563]*kernel[1]+tmp[8564]*kernel[2]+tmp[8662]*kernel[3]+tmp[8663]*kernel[4]+tmp[8664]*kernel[5]+tmp[8762]*kernel[6]+tmp[8763]*kernel[7]+tmp[8764]*kernel[8];
				ans[8664]<=tmp[8563]*kernel[0]+tmp[8564]*kernel[1]+tmp[8565]*kernel[2]+tmp[8663]*kernel[3]+tmp[8664]*kernel[4]+tmp[8665]*kernel[5]+tmp[8763]*kernel[6]+tmp[8764]*kernel[7]+tmp[8765]*kernel[8];
				ans[8665]<=tmp[8564]*kernel[0]+tmp[8565]*kernel[1]+tmp[8566]*kernel[2]+tmp[8664]*kernel[3]+tmp[8665]*kernel[4]+tmp[8666]*kernel[5]+tmp[8764]*kernel[6]+tmp[8765]*kernel[7]+tmp[8766]*kernel[8];
				ans[8666]<=tmp[8565]*kernel[0]+tmp[8566]*kernel[1]+tmp[8567]*kernel[2]+tmp[8665]*kernel[3]+tmp[8666]*kernel[4]+tmp[8667]*kernel[5]+tmp[8765]*kernel[6]+tmp[8766]*kernel[7]+tmp[8767]*kernel[8];
				ans[8667]<=tmp[8566]*kernel[0]+tmp[8567]*kernel[1]+tmp[8568]*kernel[2]+tmp[8666]*kernel[3]+tmp[8667]*kernel[4]+tmp[8668]*kernel[5]+tmp[8766]*kernel[6]+tmp[8767]*kernel[7]+tmp[8768]*kernel[8];
				ans[8668]<=tmp[8567]*kernel[0]+tmp[8568]*kernel[1]+tmp[8569]*kernel[2]+tmp[8667]*kernel[3]+tmp[8668]*kernel[4]+tmp[8669]*kernel[5]+tmp[8767]*kernel[6]+tmp[8768]*kernel[7]+tmp[8769]*kernel[8];
				ans[8669]<=tmp[8568]*kernel[0]+tmp[8569]*kernel[1]+tmp[8570]*kernel[2]+tmp[8668]*kernel[3]+tmp[8669]*kernel[4]+tmp[8670]*kernel[5]+tmp[8768]*kernel[6]+tmp[8769]*kernel[7]+tmp[8770]*kernel[8];
				ans[8670]<=tmp[8569]*kernel[0]+tmp[8570]*kernel[1]+tmp[8571]*kernel[2]+tmp[8669]*kernel[3]+tmp[8670]*kernel[4]+tmp[8671]*kernel[5]+tmp[8769]*kernel[6]+tmp[8770]*kernel[7]+tmp[8771]*kernel[8];
				ans[8671]<=tmp[8570]*kernel[0]+tmp[8571]*kernel[1]+tmp[8572]*kernel[2]+tmp[8670]*kernel[3]+tmp[8671]*kernel[4]+tmp[8672]*kernel[5]+tmp[8770]*kernel[6]+tmp[8771]*kernel[7]+tmp[8772]*kernel[8];
				ans[8672]<=tmp[8571]*kernel[0]+tmp[8572]*kernel[1]+tmp[8573]*kernel[2]+tmp[8671]*kernel[3]+tmp[8672]*kernel[4]+tmp[8673]*kernel[5]+tmp[8771]*kernel[6]+tmp[8772]*kernel[7]+tmp[8773]*kernel[8];
				ans[8673]<=tmp[8572]*kernel[0]+tmp[8573]*kernel[1]+tmp[8574]*kernel[2]+tmp[8672]*kernel[3]+tmp[8673]*kernel[4]+tmp[8674]*kernel[5]+tmp[8772]*kernel[6]+tmp[8773]*kernel[7]+tmp[8774]*kernel[8];
				ans[8674]<=tmp[8573]*kernel[0]+tmp[8574]*kernel[1]+tmp[8575]*kernel[2]+tmp[8673]*kernel[3]+tmp[8674]*kernel[4]+tmp[8675]*kernel[5]+tmp[8773]*kernel[6]+tmp[8774]*kernel[7]+tmp[8775]*kernel[8];
				ans[8675]<=tmp[8574]*kernel[0]+tmp[8575]*kernel[1]+tmp[8576]*kernel[2]+tmp[8674]*kernel[3]+tmp[8675]*kernel[4]+tmp[8676]*kernel[5]+tmp[8774]*kernel[6]+tmp[8775]*kernel[7]+tmp[8776]*kernel[8];
				ans[8676]<=tmp[8575]*kernel[0]+tmp[8576]*kernel[1]+tmp[8577]*kernel[2]+tmp[8675]*kernel[3]+tmp[8676]*kernel[4]+tmp[8677]*kernel[5]+tmp[8775]*kernel[6]+tmp[8776]*kernel[7]+tmp[8777]*kernel[8];
				ans[8677]<=tmp[8576]*kernel[0]+tmp[8577]*kernel[1]+tmp[8578]*kernel[2]+tmp[8676]*kernel[3]+tmp[8677]*kernel[4]+tmp[8678]*kernel[5]+tmp[8776]*kernel[6]+tmp[8777]*kernel[7]+tmp[8778]*kernel[8];
				ans[8678]<=tmp[8577]*kernel[0]+tmp[8578]*kernel[1]+tmp[8579]*kernel[2]+tmp[8677]*kernel[3]+tmp[8678]*kernel[4]+tmp[8679]*kernel[5]+tmp[8777]*kernel[6]+tmp[8778]*kernel[7]+tmp[8779]*kernel[8];
				ans[8679]<=tmp[8578]*kernel[0]+tmp[8579]*kernel[1]+tmp[8580]*kernel[2]+tmp[8678]*kernel[3]+tmp[8679]*kernel[4]+tmp[8680]*kernel[5]+tmp[8778]*kernel[6]+tmp[8779]*kernel[7]+tmp[8780]*kernel[8];
				ans[8680]<=tmp[8579]*kernel[0]+tmp[8580]*kernel[1]+tmp[8581]*kernel[2]+tmp[8679]*kernel[3]+tmp[8680]*kernel[4]+tmp[8681]*kernel[5]+tmp[8779]*kernel[6]+tmp[8780]*kernel[7]+tmp[8781]*kernel[8];
				ans[8681]<=tmp[8580]*kernel[0]+tmp[8581]*kernel[1]+tmp[8582]*kernel[2]+tmp[8680]*kernel[3]+tmp[8681]*kernel[4]+tmp[8682]*kernel[5]+tmp[8780]*kernel[6]+tmp[8781]*kernel[7]+tmp[8782]*kernel[8];
				ans[8682]<=tmp[8581]*kernel[0]+tmp[8582]*kernel[1]+tmp[8583]*kernel[2]+tmp[8681]*kernel[3]+tmp[8682]*kernel[4]+tmp[8683]*kernel[5]+tmp[8781]*kernel[6]+tmp[8782]*kernel[7]+tmp[8783]*kernel[8];
				ans[8683]<=tmp[8582]*kernel[0]+tmp[8583]*kernel[1]+tmp[8584]*kernel[2]+tmp[8682]*kernel[3]+tmp[8683]*kernel[4]+tmp[8684]*kernel[5]+tmp[8782]*kernel[6]+tmp[8783]*kernel[7]+tmp[8784]*kernel[8];
				ans[8684]<=tmp[8583]*kernel[0]+tmp[8584]*kernel[1]+tmp[8585]*kernel[2]+tmp[8683]*kernel[3]+tmp[8684]*kernel[4]+tmp[8685]*kernel[5]+tmp[8783]*kernel[6]+tmp[8784]*kernel[7]+tmp[8785]*kernel[8];
				ans[8685]<=tmp[8584]*kernel[0]+tmp[8585]*kernel[1]+tmp[8586]*kernel[2]+tmp[8684]*kernel[3]+tmp[8685]*kernel[4]+tmp[8686]*kernel[5]+tmp[8784]*kernel[6]+tmp[8785]*kernel[7]+tmp[8786]*kernel[8];
				ans[8686]<=tmp[8585]*kernel[0]+tmp[8586]*kernel[1]+tmp[8587]*kernel[2]+tmp[8685]*kernel[3]+tmp[8686]*kernel[4]+tmp[8687]*kernel[5]+tmp[8785]*kernel[6]+tmp[8786]*kernel[7]+tmp[8787]*kernel[8];
				ans[8687]<=tmp[8586]*kernel[0]+tmp[8587]*kernel[1]+tmp[8588]*kernel[2]+tmp[8686]*kernel[3]+tmp[8687]*kernel[4]+tmp[8688]*kernel[5]+tmp[8786]*kernel[6]+tmp[8787]*kernel[7]+tmp[8788]*kernel[8];
				ans[8688]<=tmp[8587]*kernel[0]+tmp[8588]*kernel[1]+tmp[8589]*kernel[2]+tmp[8687]*kernel[3]+tmp[8688]*kernel[4]+tmp[8689]*kernel[5]+tmp[8787]*kernel[6]+tmp[8788]*kernel[7]+tmp[8789]*kernel[8];
				ans[8689]<=tmp[8588]*kernel[0]+tmp[8589]*kernel[1]+tmp[8590]*kernel[2]+tmp[8688]*kernel[3]+tmp[8689]*kernel[4]+tmp[8690]*kernel[5]+tmp[8788]*kernel[6]+tmp[8789]*kernel[7]+tmp[8790]*kernel[8];
				ans[8690]<=tmp[8589]*kernel[0]+tmp[8590]*kernel[1]+tmp[8591]*kernel[2]+tmp[8689]*kernel[3]+tmp[8690]*kernel[4]+tmp[8691]*kernel[5]+tmp[8789]*kernel[6]+tmp[8790]*kernel[7]+tmp[8791]*kernel[8];
				ans[8691]<=tmp[8590]*kernel[0]+tmp[8591]*kernel[1]+tmp[8592]*kernel[2]+tmp[8690]*kernel[3]+tmp[8691]*kernel[4]+tmp[8692]*kernel[5]+tmp[8790]*kernel[6]+tmp[8791]*kernel[7]+tmp[8792]*kernel[8];
				ans[8692]<=tmp[8591]*kernel[0]+tmp[8592]*kernel[1]+tmp[8593]*kernel[2]+tmp[8691]*kernel[3]+tmp[8692]*kernel[4]+tmp[8693]*kernel[5]+tmp[8791]*kernel[6]+tmp[8792]*kernel[7]+tmp[8793]*kernel[8];
				ans[8693]<=tmp[8592]*kernel[0]+tmp[8593]*kernel[1]+tmp[8594]*kernel[2]+tmp[8692]*kernel[3]+tmp[8693]*kernel[4]+tmp[8694]*kernel[5]+tmp[8792]*kernel[6]+tmp[8793]*kernel[7]+tmp[8794]*kernel[8];
				ans[8694]<=tmp[8593]*kernel[0]+tmp[8594]*kernel[1]+tmp[8595]*kernel[2]+tmp[8693]*kernel[3]+tmp[8694]*kernel[4]+tmp[8695]*kernel[5]+tmp[8793]*kernel[6]+tmp[8794]*kernel[7]+tmp[8795]*kernel[8];
				ans[8695]<=tmp[8594]*kernel[0]+tmp[8595]*kernel[1]+tmp[8596]*kernel[2]+tmp[8694]*kernel[3]+tmp[8695]*kernel[4]+tmp[8696]*kernel[5]+tmp[8794]*kernel[6]+tmp[8795]*kernel[7]+tmp[8796]*kernel[8];
				ans[8696]<=tmp[8595]*kernel[0]+tmp[8596]*kernel[1]+tmp[8597]*kernel[2]+tmp[8695]*kernel[3]+tmp[8696]*kernel[4]+tmp[8697]*kernel[5]+tmp[8795]*kernel[6]+tmp[8796]*kernel[7]+tmp[8797]*kernel[8];
				ans[8697]<=tmp[8596]*kernel[0]+tmp[8597]*kernel[1]+tmp[8598]*kernel[2]+tmp[8696]*kernel[3]+tmp[8697]*kernel[4]+tmp[8698]*kernel[5]+tmp[8796]*kernel[6]+tmp[8797]*kernel[7]+tmp[8798]*kernel[8];
				ans[8698]<=tmp[8597]*kernel[0]+tmp[8598]*kernel[1]+tmp[8599]*kernel[2]+tmp[8697]*kernel[3]+tmp[8698]*kernel[4]+tmp[8699]*kernel[5]+tmp[8797]*kernel[6]+tmp[8798]*kernel[7]+tmp[8799]*kernel[8];
				ans[8699]<=tmp[8598]*kernel[0]+tmp[8599]*kernel[1]+tmp[8698]*kernel[3]+tmp[8699]*kernel[4]+tmp[8798]*kernel[6]+tmp[8799]*kernel[7];
				ans[8700]<=tmp[8600]*kernel[1]+tmp[8601]*kernel[2]+tmp[8700]*kernel[4]+tmp[8701]*kernel[5]+tmp[8800]*kernel[7]+tmp[8801]*kernel[8];
				ans[8701]<=tmp[8600]*kernel[0]+tmp[8601]*kernel[1]+tmp[8602]*kernel[2]+tmp[8700]*kernel[3]+tmp[8701]*kernel[4]+tmp[8702]*kernel[5]+tmp[8800]*kernel[6]+tmp[8801]*kernel[7]+tmp[8802]*kernel[8];
				ans[8702]<=tmp[8601]*kernel[0]+tmp[8602]*kernel[1]+tmp[8603]*kernel[2]+tmp[8701]*kernel[3]+tmp[8702]*kernel[4]+tmp[8703]*kernel[5]+tmp[8801]*kernel[6]+tmp[8802]*kernel[7]+tmp[8803]*kernel[8];
				ans[8703]<=tmp[8602]*kernel[0]+tmp[8603]*kernel[1]+tmp[8604]*kernel[2]+tmp[8702]*kernel[3]+tmp[8703]*kernel[4]+tmp[8704]*kernel[5]+tmp[8802]*kernel[6]+tmp[8803]*kernel[7]+tmp[8804]*kernel[8];
				ans[8704]<=tmp[8603]*kernel[0]+tmp[8604]*kernel[1]+tmp[8605]*kernel[2]+tmp[8703]*kernel[3]+tmp[8704]*kernel[4]+tmp[8705]*kernel[5]+tmp[8803]*kernel[6]+tmp[8804]*kernel[7]+tmp[8805]*kernel[8];
				ans[8705]<=tmp[8604]*kernel[0]+tmp[8605]*kernel[1]+tmp[8606]*kernel[2]+tmp[8704]*kernel[3]+tmp[8705]*kernel[4]+tmp[8706]*kernel[5]+tmp[8804]*kernel[6]+tmp[8805]*kernel[7]+tmp[8806]*kernel[8];
				ans[8706]<=tmp[8605]*kernel[0]+tmp[8606]*kernel[1]+tmp[8607]*kernel[2]+tmp[8705]*kernel[3]+tmp[8706]*kernel[4]+tmp[8707]*kernel[5]+tmp[8805]*kernel[6]+tmp[8806]*kernel[7]+tmp[8807]*kernel[8];
				ans[8707]<=tmp[8606]*kernel[0]+tmp[8607]*kernel[1]+tmp[8608]*kernel[2]+tmp[8706]*kernel[3]+tmp[8707]*kernel[4]+tmp[8708]*kernel[5]+tmp[8806]*kernel[6]+tmp[8807]*kernel[7]+tmp[8808]*kernel[8];
				ans[8708]<=tmp[8607]*kernel[0]+tmp[8608]*kernel[1]+tmp[8609]*kernel[2]+tmp[8707]*kernel[3]+tmp[8708]*kernel[4]+tmp[8709]*kernel[5]+tmp[8807]*kernel[6]+tmp[8808]*kernel[7]+tmp[8809]*kernel[8];
				ans[8709]<=tmp[8608]*kernel[0]+tmp[8609]*kernel[1]+tmp[8610]*kernel[2]+tmp[8708]*kernel[3]+tmp[8709]*kernel[4]+tmp[8710]*kernel[5]+tmp[8808]*kernel[6]+tmp[8809]*kernel[7]+tmp[8810]*kernel[8];
				ans[8710]<=tmp[8609]*kernel[0]+tmp[8610]*kernel[1]+tmp[8611]*kernel[2]+tmp[8709]*kernel[3]+tmp[8710]*kernel[4]+tmp[8711]*kernel[5]+tmp[8809]*kernel[6]+tmp[8810]*kernel[7]+tmp[8811]*kernel[8];
				ans[8711]<=tmp[8610]*kernel[0]+tmp[8611]*kernel[1]+tmp[8612]*kernel[2]+tmp[8710]*kernel[3]+tmp[8711]*kernel[4]+tmp[8712]*kernel[5]+tmp[8810]*kernel[6]+tmp[8811]*kernel[7]+tmp[8812]*kernel[8];
				ans[8712]<=tmp[8611]*kernel[0]+tmp[8612]*kernel[1]+tmp[8613]*kernel[2]+tmp[8711]*kernel[3]+tmp[8712]*kernel[4]+tmp[8713]*kernel[5]+tmp[8811]*kernel[6]+tmp[8812]*kernel[7]+tmp[8813]*kernel[8];
				ans[8713]<=tmp[8612]*kernel[0]+tmp[8613]*kernel[1]+tmp[8614]*kernel[2]+tmp[8712]*kernel[3]+tmp[8713]*kernel[4]+tmp[8714]*kernel[5]+tmp[8812]*kernel[6]+tmp[8813]*kernel[7]+tmp[8814]*kernel[8];
				ans[8714]<=tmp[8613]*kernel[0]+tmp[8614]*kernel[1]+tmp[8615]*kernel[2]+tmp[8713]*kernel[3]+tmp[8714]*kernel[4]+tmp[8715]*kernel[5]+tmp[8813]*kernel[6]+tmp[8814]*kernel[7]+tmp[8815]*kernel[8];
				ans[8715]<=tmp[8614]*kernel[0]+tmp[8615]*kernel[1]+tmp[8616]*kernel[2]+tmp[8714]*kernel[3]+tmp[8715]*kernel[4]+tmp[8716]*kernel[5]+tmp[8814]*kernel[6]+tmp[8815]*kernel[7]+tmp[8816]*kernel[8];
				ans[8716]<=tmp[8615]*kernel[0]+tmp[8616]*kernel[1]+tmp[8617]*kernel[2]+tmp[8715]*kernel[3]+tmp[8716]*kernel[4]+tmp[8717]*kernel[5]+tmp[8815]*kernel[6]+tmp[8816]*kernel[7]+tmp[8817]*kernel[8];
				ans[8717]<=tmp[8616]*kernel[0]+tmp[8617]*kernel[1]+tmp[8618]*kernel[2]+tmp[8716]*kernel[3]+tmp[8717]*kernel[4]+tmp[8718]*kernel[5]+tmp[8816]*kernel[6]+tmp[8817]*kernel[7]+tmp[8818]*kernel[8];
				ans[8718]<=tmp[8617]*kernel[0]+tmp[8618]*kernel[1]+tmp[8619]*kernel[2]+tmp[8717]*kernel[3]+tmp[8718]*kernel[4]+tmp[8719]*kernel[5]+tmp[8817]*kernel[6]+tmp[8818]*kernel[7]+tmp[8819]*kernel[8];
				ans[8719]<=tmp[8618]*kernel[0]+tmp[8619]*kernel[1]+tmp[8620]*kernel[2]+tmp[8718]*kernel[3]+tmp[8719]*kernel[4]+tmp[8720]*kernel[5]+tmp[8818]*kernel[6]+tmp[8819]*kernel[7]+tmp[8820]*kernel[8];
				ans[8720]<=tmp[8619]*kernel[0]+tmp[8620]*kernel[1]+tmp[8621]*kernel[2]+tmp[8719]*kernel[3]+tmp[8720]*kernel[4]+tmp[8721]*kernel[5]+tmp[8819]*kernel[6]+tmp[8820]*kernel[7]+tmp[8821]*kernel[8];
				ans[8721]<=tmp[8620]*kernel[0]+tmp[8621]*kernel[1]+tmp[8622]*kernel[2]+tmp[8720]*kernel[3]+tmp[8721]*kernel[4]+tmp[8722]*kernel[5]+tmp[8820]*kernel[6]+tmp[8821]*kernel[7]+tmp[8822]*kernel[8];
				ans[8722]<=tmp[8621]*kernel[0]+tmp[8622]*kernel[1]+tmp[8623]*kernel[2]+tmp[8721]*kernel[3]+tmp[8722]*kernel[4]+tmp[8723]*kernel[5]+tmp[8821]*kernel[6]+tmp[8822]*kernel[7]+tmp[8823]*kernel[8];
				ans[8723]<=tmp[8622]*kernel[0]+tmp[8623]*kernel[1]+tmp[8624]*kernel[2]+tmp[8722]*kernel[3]+tmp[8723]*kernel[4]+tmp[8724]*kernel[5]+tmp[8822]*kernel[6]+tmp[8823]*kernel[7]+tmp[8824]*kernel[8];
				ans[8724]<=tmp[8623]*kernel[0]+tmp[8624]*kernel[1]+tmp[8625]*kernel[2]+tmp[8723]*kernel[3]+tmp[8724]*kernel[4]+tmp[8725]*kernel[5]+tmp[8823]*kernel[6]+tmp[8824]*kernel[7]+tmp[8825]*kernel[8];
				ans[8725]<=tmp[8624]*kernel[0]+tmp[8625]*kernel[1]+tmp[8626]*kernel[2]+tmp[8724]*kernel[3]+tmp[8725]*kernel[4]+tmp[8726]*kernel[5]+tmp[8824]*kernel[6]+tmp[8825]*kernel[7]+tmp[8826]*kernel[8];
				ans[8726]<=tmp[8625]*kernel[0]+tmp[8626]*kernel[1]+tmp[8627]*kernel[2]+tmp[8725]*kernel[3]+tmp[8726]*kernel[4]+tmp[8727]*kernel[5]+tmp[8825]*kernel[6]+tmp[8826]*kernel[7]+tmp[8827]*kernel[8];
				ans[8727]<=tmp[8626]*kernel[0]+tmp[8627]*kernel[1]+tmp[8628]*kernel[2]+tmp[8726]*kernel[3]+tmp[8727]*kernel[4]+tmp[8728]*kernel[5]+tmp[8826]*kernel[6]+tmp[8827]*kernel[7]+tmp[8828]*kernel[8];
				ans[8728]<=tmp[8627]*kernel[0]+tmp[8628]*kernel[1]+tmp[8629]*kernel[2]+tmp[8727]*kernel[3]+tmp[8728]*kernel[4]+tmp[8729]*kernel[5]+tmp[8827]*kernel[6]+tmp[8828]*kernel[7]+tmp[8829]*kernel[8];
				ans[8729]<=tmp[8628]*kernel[0]+tmp[8629]*kernel[1]+tmp[8630]*kernel[2]+tmp[8728]*kernel[3]+tmp[8729]*kernel[4]+tmp[8730]*kernel[5]+tmp[8828]*kernel[6]+tmp[8829]*kernel[7]+tmp[8830]*kernel[8];
				ans[8730]<=tmp[8629]*kernel[0]+tmp[8630]*kernel[1]+tmp[8631]*kernel[2]+tmp[8729]*kernel[3]+tmp[8730]*kernel[4]+tmp[8731]*kernel[5]+tmp[8829]*kernel[6]+tmp[8830]*kernel[7]+tmp[8831]*kernel[8];
				ans[8731]<=tmp[8630]*kernel[0]+tmp[8631]*kernel[1]+tmp[8632]*kernel[2]+tmp[8730]*kernel[3]+tmp[8731]*kernel[4]+tmp[8732]*kernel[5]+tmp[8830]*kernel[6]+tmp[8831]*kernel[7]+tmp[8832]*kernel[8];
				ans[8732]<=tmp[8631]*kernel[0]+tmp[8632]*kernel[1]+tmp[8633]*kernel[2]+tmp[8731]*kernel[3]+tmp[8732]*kernel[4]+tmp[8733]*kernel[5]+tmp[8831]*kernel[6]+tmp[8832]*kernel[7]+tmp[8833]*kernel[8];
				ans[8733]<=tmp[8632]*kernel[0]+tmp[8633]*kernel[1]+tmp[8634]*kernel[2]+tmp[8732]*kernel[3]+tmp[8733]*kernel[4]+tmp[8734]*kernel[5]+tmp[8832]*kernel[6]+tmp[8833]*kernel[7]+tmp[8834]*kernel[8];
				ans[8734]<=tmp[8633]*kernel[0]+tmp[8634]*kernel[1]+tmp[8635]*kernel[2]+tmp[8733]*kernel[3]+tmp[8734]*kernel[4]+tmp[8735]*kernel[5]+tmp[8833]*kernel[6]+tmp[8834]*kernel[7]+tmp[8835]*kernel[8];
				ans[8735]<=tmp[8634]*kernel[0]+tmp[8635]*kernel[1]+tmp[8636]*kernel[2]+tmp[8734]*kernel[3]+tmp[8735]*kernel[4]+tmp[8736]*kernel[5]+tmp[8834]*kernel[6]+tmp[8835]*kernel[7]+tmp[8836]*kernel[8];
				ans[8736]<=tmp[8635]*kernel[0]+tmp[8636]*kernel[1]+tmp[8637]*kernel[2]+tmp[8735]*kernel[3]+tmp[8736]*kernel[4]+tmp[8737]*kernel[5]+tmp[8835]*kernel[6]+tmp[8836]*kernel[7]+tmp[8837]*kernel[8];
				ans[8737]<=tmp[8636]*kernel[0]+tmp[8637]*kernel[1]+tmp[8638]*kernel[2]+tmp[8736]*kernel[3]+tmp[8737]*kernel[4]+tmp[8738]*kernel[5]+tmp[8836]*kernel[6]+tmp[8837]*kernel[7]+tmp[8838]*kernel[8];
				ans[8738]<=tmp[8637]*kernel[0]+tmp[8638]*kernel[1]+tmp[8639]*kernel[2]+tmp[8737]*kernel[3]+tmp[8738]*kernel[4]+tmp[8739]*kernel[5]+tmp[8837]*kernel[6]+tmp[8838]*kernel[7]+tmp[8839]*kernel[8];
				ans[8739]<=tmp[8638]*kernel[0]+tmp[8639]*kernel[1]+tmp[8640]*kernel[2]+tmp[8738]*kernel[3]+tmp[8739]*kernel[4]+tmp[8740]*kernel[5]+tmp[8838]*kernel[6]+tmp[8839]*kernel[7]+tmp[8840]*kernel[8];
				ans[8740]<=tmp[8639]*kernel[0]+tmp[8640]*kernel[1]+tmp[8641]*kernel[2]+tmp[8739]*kernel[3]+tmp[8740]*kernel[4]+tmp[8741]*kernel[5]+tmp[8839]*kernel[6]+tmp[8840]*kernel[7]+tmp[8841]*kernel[8];
				ans[8741]<=tmp[8640]*kernel[0]+tmp[8641]*kernel[1]+tmp[8642]*kernel[2]+tmp[8740]*kernel[3]+tmp[8741]*kernel[4]+tmp[8742]*kernel[5]+tmp[8840]*kernel[6]+tmp[8841]*kernel[7]+tmp[8842]*kernel[8];
				ans[8742]<=tmp[8641]*kernel[0]+tmp[8642]*kernel[1]+tmp[8643]*kernel[2]+tmp[8741]*kernel[3]+tmp[8742]*kernel[4]+tmp[8743]*kernel[5]+tmp[8841]*kernel[6]+tmp[8842]*kernel[7]+tmp[8843]*kernel[8];
				ans[8743]<=tmp[8642]*kernel[0]+tmp[8643]*kernel[1]+tmp[8644]*kernel[2]+tmp[8742]*kernel[3]+tmp[8743]*kernel[4]+tmp[8744]*kernel[5]+tmp[8842]*kernel[6]+tmp[8843]*kernel[7]+tmp[8844]*kernel[8];
				ans[8744]<=tmp[8643]*kernel[0]+tmp[8644]*kernel[1]+tmp[8645]*kernel[2]+tmp[8743]*kernel[3]+tmp[8744]*kernel[4]+tmp[8745]*kernel[5]+tmp[8843]*kernel[6]+tmp[8844]*kernel[7]+tmp[8845]*kernel[8];
				ans[8745]<=tmp[8644]*kernel[0]+tmp[8645]*kernel[1]+tmp[8646]*kernel[2]+tmp[8744]*kernel[3]+tmp[8745]*kernel[4]+tmp[8746]*kernel[5]+tmp[8844]*kernel[6]+tmp[8845]*kernel[7]+tmp[8846]*kernel[8];
				ans[8746]<=tmp[8645]*kernel[0]+tmp[8646]*kernel[1]+tmp[8647]*kernel[2]+tmp[8745]*kernel[3]+tmp[8746]*kernel[4]+tmp[8747]*kernel[5]+tmp[8845]*kernel[6]+tmp[8846]*kernel[7]+tmp[8847]*kernel[8];
				ans[8747]<=tmp[8646]*kernel[0]+tmp[8647]*kernel[1]+tmp[8648]*kernel[2]+tmp[8746]*kernel[3]+tmp[8747]*kernel[4]+tmp[8748]*kernel[5]+tmp[8846]*kernel[6]+tmp[8847]*kernel[7]+tmp[8848]*kernel[8];
				ans[8748]<=tmp[8647]*kernel[0]+tmp[8648]*kernel[1]+tmp[8649]*kernel[2]+tmp[8747]*kernel[3]+tmp[8748]*kernel[4]+tmp[8749]*kernel[5]+tmp[8847]*kernel[6]+tmp[8848]*kernel[7]+tmp[8849]*kernel[8];
				ans[8749]<=tmp[8648]*kernel[0]+tmp[8649]*kernel[1]+tmp[8650]*kernel[2]+tmp[8748]*kernel[3]+tmp[8749]*kernel[4]+tmp[8750]*kernel[5]+tmp[8848]*kernel[6]+tmp[8849]*kernel[7]+tmp[8850]*kernel[8];
				ans[8750]<=tmp[8649]*kernel[0]+tmp[8650]*kernel[1]+tmp[8651]*kernel[2]+tmp[8749]*kernel[3]+tmp[8750]*kernel[4]+tmp[8751]*kernel[5]+tmp[8849]*kernel[6]+tmp[8850]*kernel[7]+tmp[8851]*kernel[8];
				ans[8751]<=tmp[8650]*kernel[0]+tmp[8651]*kernel[1]+tmp[8652]*kernel[2]+tmp[8750]*kernel[3]+tmp[8751]*kernel[4]+tmp[8752]*kernel[5]+tmp[8850]*kernel[6]+tmp[8851]*kernel[7]+tmp[8852]*kernel[8];
				ans[8752]<=tmp[8651]*kernel[0]+tmp[8652]*kernel[1]+tmp[8653]*kernel[2]+tmp[8751]*kernel[3]+tmp[8752]*kernel[4]+tmp[8753]*kernel[5]+tmp[8851]*kernel[6]+tmp[8852]*kernel[7]+tmp[8853]*kernel[8];
				ans[8753]<=tmp[8652]*kernel[0]+tmp[8653]*kernel[1]+tmp[8654]*kernel[2]+tmp[8752]*kernel[3]+tmp[8753]*kernel[4]+tmp[8754]*kernel[5]+tmp[8852]*kernel[6]+tmp[8853]*kernel[7]+tmp[8854]*kernel[8];
				ans[8754]<=tmp[8653]*kernel[0]+tmp[8654]*kernel[1]+tmp[8655]*kernel[2]+tmp[8753]*kernel[3]+tmp[8754]*kernel[4]+tmp[8755]*kernel[5]+tmp[8853]*kernel[6]+tmp[8854]*kernel[7]+tmp[8855]*kernel[8];
				ans[8755]<=tmp[8654]*kernel[0]+tmp[8655]*kernel[1]+tmp[8656]*kernel[2]+tmp[8754]*kernel[3]+tmp[8755]*kernel[4]+tmp[8756]*kernel[5]+tmp[8854]*kernel[6]+tmp[8855]*kernel[7]+tmp[8856]*kernel[8];
				ans[8756]<=tmp[8655]*kernel[0]+tmp[8656]*kernel[1]+tmp[8657]*kernel[2]+tmp[8755]*kernel[3]+tmp[8756]*kernel[4]+tmp[8757]*kernel[5]+tmp[8855]*kernel[6]+tmp[8856]*kernel[7]+tmp[8857]*kernel[8];
				ans[8757]<=tmp[8656]*kernel[0]+tmp[8657]*kernel[1]+tmp[8658]*kernel[2]+tmp[8756]*kernel[3]+tmp[8757]*kernel[4]+tmp[8758]*kernel[5]+tmp[8856]*kernel[6]+tmp[8857]*kernel[7]+tmp[8858]*kernel[8];
				ans[8758]<=tmp[8657]*kernel[0]+tmp[8658]*kernel[1]+tmp[8659]*kernel[2]+tmp[8757]*kernel[3]+tmp[8758]*kernel[4]+tmp[8759]*kernel[5]+tmp[8857]*kernel[6]+tmp[8858]*kernel[7]+tmp[8859]*kernel[8];
				ans[8759]<=tmp[8658]*kernel[0]+tmp[8659]*kernel[1]+tmp[8660]*kernel[2]+tmp[8758]*kernel[3]+tmp[8759]*kernel[4]+tmp[8760]*kernel[5]+tmp[8858]*kernel[6]+tmp[8859]*kernel[7]+tmp[8860]*kernel[8];
				ans[8760]<=tmp[8659]*kernel[0]+tmp[8660]*kernel[1]+tmp[8661]*kernel[2]+tmp[8759]*kernel[3]+tmp[8760]*kernel[4]+tmp[8761]*kernel[5]+tmp[8859]*kernel[6]+tmp[8860]*kernel[7]+tmp[8861]*kernel[8];
				ans[8761]<=tmp[8660]*kernel[0]+tmp[8661]*kernel[1]+tmp[8662]*kernel[2]+tmp[8760]*kernel[3]+tmp[8761]*kernel[4]+tmp[8762]*kernel[5]+tmp[8860]*kernel[6]+tmp[8861]*kernel[7]+tmp[8862]*kernel[8];
				ans[8762]<=tmp[8661]*kernel[0]+tmp[8662]*kernel[1]+tmp[8663]*kernel[2]+tmp[8761]*kernel[3]+tmp[8762]*kernel[4]+tmp[8763]*kernel[5]+tmp[8861]*kernel[6]+tmp[8862]*kernel[7]+tmp[8863]*kernel[8];
				ans[8763]<=tmp[8662]*kernel[0]+tmp[8663]*kernel[1]+tmp[8664]*kernel[2]+tmp[8762]*kernel[3]+tmp[8763]*kernel[4]+tmp[8764]*kernel[5]+tmp[8862]*kernel[6]+tmp[8863]*kernel[7]+tmp[8864]*kernel[8];
				ans[8764]<=tmp[8663]*kernel[0]+tmp[8664]*kernel[1]+tmp[8665]*kernel[2]+tmp[8763]*kernel[3]+tmp[8764]*kernel[4]+tmp[8765]*kernel[5]+tmp[8863]*kernel[6]+tmp[8864]*kernel[7]+tmp[8865]*kernel[8];
				ans[8765]<=tmp[8664]*kernel[0]+tmp[8665]*kernel[1]+tmp[8666]*kernel[2]+tmp[8764]*kernel[3]+tmp[8765]*kernel[4]+tmp[8766]*kernel[5]+tmp[8864]*kernel[6]+tmp[8865]*kernel[7]+tmp[8866]*kernel[8];
				ans[8766]<=tmp[8665]*kernel[0]+tmp[8666]*kernel[1]+tmp[8667]*kernel[2]+tmp[8765]*kernel[3]+tmp[8766]*kernel[4]+tmp[8767]*kernel[5]+tmp[8865]*kernel[6]+tmp[8866]*kernel[7]+tmp[8867]*kernel[8];
				ans[8767]<=tmp[8666]*kernel[0]+tmp[8667]*kernel[1]+tmp[8668]*kernel[2]+tmp[8766]*kernel[3]+tmp[8767]*kernel[4]+tmp[8768]*kernel[5]+tmp[8866]*kernel[6]+tmp[8867]*kernel[7]+tmp[8868]*kernel[8];
				ans[8768]<=tmp[8667]*kernel[0]+tmp[8668]*kernel[1]+tmp[8669]*kernel[2]+tmp[8767]*kernel[3]+tmp[8768]*kernel[4]+tmp[8769]*kernel[5]+tmp[8867]*kernel[6]+tmp[8868]*kernel[7]+tmp[8869]*kernel[8];
				ans[8769]<=tmp[8668]*kernel[0]+tmp[8669]*kernel[1]+tmp[8670]*kernel[2]+tmp[8768]*kernel[3]+tmp[8769]*kernel[4]+tmp[8770]*kernel[5]+tmp[8868]*kernel[6]+tmp[8869]*kernel[7]+tmp[8870]*kernel[8];
				ans[8770]<=tmp[8669]*kernel[0]+tmp[8670]*kernel[1]+tmp[8671]*kernel[2]+tmp[8769]*kernel[3]+tmp[8770]*kernel[4]+tmp[8771]*kernel[5]+tmp[8869]*kernel[6]+tmp[8870]*kernel[7]+tmp[8871]*kernel[8];
				ans[8771]<=tmp[8670]*kernel[0]+tmp[8671]*kernel[1]+tmp[8672]*kernel[2]+tmp[8770]*kernel[3]+tmp[8771]*kernel[4]+tmp[8772]*kernel[5]+tmp[8870]*kernel[6]+tmp[8871]*kernel[7]+tmp[8872]*kernel[8];
				ans[8772]<=tmp[8671]*kernel[0]+tmp[8672]*kernel[1]+tmp[8673]*kernel[2]+tmp[8771]*kernel[3]+tmp[8772]*kernel[4]+tmp[8773]*kernel[5]+tmp[8871]*kernel[6]+tmp[8872]*kernel[7]+tmp[8873]*kernel[8];
				ans[8773]<=tmp[8672]*kernel[0]+tmp[8673]*kernel[1]+tmp[8674]*kernel[2]+tmp[8772]*kernel[3]+tmp[8773]*kernel[4]+tmp[8774]*kernel[5]+tmp[8872]*kernel[6]+tmp[8873]*kernel[7]+tmp[8874]*kernel[8];
				ans[8774]<=tmp[8673]*kernel[0]+tmp[8674]*kernel[1]+tmp[8675]*kernel[2]+tmp[8773]*kernel[3]+tmp[8774]*kernel[4]+tmp[8775]*kernel[5]+tmp[8873]*kernel[6]+tmp[8874]*kernel[7]+tmp[8875]*kernel[8];
				ans[8775]<=tmp[8674]*kernel[0]+tmp[8675]*kernel[1]+tmp[8676]*kernel[2]+tmp[8774]*kernel[3]+tmp[8775]*kernel[4]+tmp[8776]*kernel[5]+tmp[8874]*kernel[6]+tmp[8875]*kernel[7]+tmp[8876]*kernel[8];
				ans[8776]<=tmp[8675]*kernel[0]+tmp[8676]*kernel[1]+tmp[8677]*kernel[2]+tmp[8775]*kernel[3]+tmp[8776]*kernel[4]+tmp[8777]*kernel[5]+tmp[8875]*kernel[6]+tmp[8876]*kernel[7]+tmp[8877]*kernel[8];
				ans[8777]<=tmp[8676]*kernel[0]+tmp[8677]*kernel[1]+tmp[8678]*kernel[2]+tmp[8776]*kernel[3]+tmp[8777]*kernel[4]+tmp[8778]*kernel[5]+tmp[8876]*kernel[6]+tmp[8877]*kernel[7]+tmp[8878]*kernel[8];
				ans[8778]<=tmp[8677]*kernel[0]+tmp[8678]*kernel[1]+tmp[8679]*kernel[2]+tmp[8777]*kernel[3]+tmp[8778]*kernel[4]+tmp[8779]*kernel[5]+tmp[8877]*kernel[6]+tmp[8878]*kernel[7]+tmp[8879]*kernel[8];
				ans[8779]<=tmp[8678]*kernel[0]+tmp[8679]*kernel[1]+tmp[8680]*kernel[2]+tmp[8778]*kernel[3]+tmp[8779]*kernel[4]+tmp[8780]*kernel[5]+tmp[8878]*kernel[6]+tmp[8879]*kernel[7]+tmp[8880]*kernel[8];
				ans[8780]<=tmp[8679]*kernel[0]+tmp[8680]*kernel[1]+tmp[8681]*kernel[2]+tmp[8779]*kernel[3]+tmp[8780]*kernel[4]+tmp[8781]*kernel[5]+tmp[8879]*kernel[6]+tmp[8880]*kernel[7]+tmp[8881]*kernel[8];
				ans[8781]<=tmp[8680]*kernel[0]+tmp[8681]*kernel[1]+tmp[8682]*kernel[2]+tmp[8780]*kernel[3]+tmp[8781]*kernel[4]+tmp[8782]*kernel[5]+tmp[8880]*kernel[6]+tmp[8881]*kernel[7]+tmp[8882]*kernel[8];
				ans[8782]<=tmp[8681]*kernel[0]+tmp[8682]*kernel[1]+tmp[8683]*kernel[2]+tmp[8781]*kernel[3]+tmp[8782]*kernel[4]+tmp[8783]*kernel[5]+tmp[8881]*kernel[6]+tmp[8882]*kernel[7]+tmp[8883]*kernel[8];
				ans[8783]<=tmp[8682]*kernel[0]+tmp[8683]*kernel[1]+tmp[8684]*kernel[2]+tmp[8782]*kernel[3]+tmp[8783]*kernel[4]+tmp[8784]*kernel[5]+tmp[8882]*kernel[6]+tmp[8883]*kernel[7]+tmp[8884]*kernel[8];
				ans[8784]<=tmp[8683]*kernel[0]+tmp[8684]*kernel[1]+tmp[8685]*kernel[2]+tmp[8783]*kernel[3]+tmp[8784]*kernel[4]+tmp[8785]*kernel[5]+tmp[8883]*kernel[6]+tmp[8884]*kernel[7]+tmp[8885]*kernel[8];
				ans[8785]<=tmp[8684]*kernel[0]+tmp[8685]*kernel[1]+tmp[8686]*kernel[2]+tmp[8784]*kernel[3]+tmp[8785]*kernel[4]+tmp[8786]*kernel[5]+tmp[8884]*kernel[6]+tmp[8885]*kernel[7]+tmp[8886]*kernel[8];
				ans[8786]<=tmp[8685]*kernel[0]+tmp[8686]*kernel[1]+tmp[8687]*kernel[2]+tmp[8785]*kernel[3]+tmp[8786]*kernel[4]+tmp[8787]*kernel[5]+tmp[8885]*kernel[6]+tmp[8886]*kernel[7]+tmp[8887]*kernel[8];
				ans[8787]<=tmp[8686]*kernel[0]+tmp[8687]*kernel[1]+tmp[8688]*kernel[2]+tmp[8786]*kernel[3]+tmp[8787]*kernel[4]+tmp[8788]*kernel[5]+tmp[8886]*kernel[6]+tmp[8887]*kernel[7]+tmp[8888]*kernel[8];
				ans[8788]<=tmp[8687]*kernel[0]+tmp[8688]*kernel[1]+tmp[8689]*kernel[2]+tmp[8787]*kernel[3]+tmp[8788]*kernel[4]+tmp[8789]*kernel[5]+tmp[8887]*kernel[6]+tmp[8888]*kernel[7]+tmp[8889]*kernel[8];
				ans[8789]<=tmp[8688]*kernel[0]+tmp[8689]*kernel[1]+tmp[8690]*kernel[2]+tmp[8788]*kernel[3]+tmp[8789]*kernel[4]+tmp[8790]*kernel[5]+tmp[8888]*kernel[6]+tmp[8889]*kernel[7]+tmp[8890]*kernel[8];
				ans[8790]<=tmp[8689]*kernel[0]+tmp[8690]*kernel[1]+tmp[8691]*kernel[2]+tmp[8789]*kernel[3]+tmp[8790]*kernel[4]+tmp[8791]*kernel[5]+tmp[8889]*kernel[6]+tmp[8890]*kernel[7]+tmp[8891]*kernel[8];
				ans[8791]<=tmp[8690]*kernel[0]+tmp[8691]*kernel[1]+tmp[8692]*kernel[2]+tmp[8790]*kernel[3]+tmp[8791]*kernel[4]+tmp[8792]*kernel[5]+tmp[8890]*kernel[6]+tmp[8891]*kernel[7]+tmp[8892]*kernel[8];
				ans[8792]<=tmp[8691]*kernel[0]+tmp[8692]*kernel[1]+tmp[8693]*kernel[2]+tmp[8791]*kernel[3]+tmp[8792]*kernel[4]+tmp[8793]*kernel[5]+tmp[8891]*kernel[6]+tmp[8892]*kernel[7]+tmp[8893]*kernel[8];
				ans[8793]<=tmp[8692]*kernel[0]+tmp[8693]*kernel[1]+tmp[8694]*kernel[2]+tmp[8792]*kernel[3]+tmp[8793]*kernel[4]+tmp[8794]*kernel[5]+tmp[8892]*kernel[6]+tmp[8893]*kernel[7]+tmp[8894]*kernel[8];
				ans[8794]<=tmp[8693]*kernel[0]+tmp[8694]*kernel[1]+tmp[8695]*kernel[2]+tmp[8793]*kernel[3]+tmp[8794]*kernel[4]+tmp[8795]*kernel[5]+tmp[8893]*kernel[6]+tmp[8894]*kernel[7]+tmp[8895]*kernel[8];
				ans[8795]<=tmp[8694]*kernel[0]+tmp[8695]*kernel[1]+tmp[8696]*kernel[2]+tmp[8794]*kernel[3]+tmp[8795]*kernel[4]+tmp[8796]*kernel[5]+tmp[8894]*kernel[6]+tmp[8895]*kernel[7]+tmp[8896]*kernel[8];
				ans[8796]<=tmp[8695]*kernel[0]+tmp[8696]*kernel[1]+tmp[8697]*kernel[2]+tmp[8795]*kernel[3]+tmp[8796]*kernel[4]+tmp[8797]*kernel[5]+tmp[8895]*kernel[6]+tmp[8896]*kernel[7]+tmp[8897]*kernel[8];
				ans[8797]<=tmp[8696]*kernel[0]+tmp[8697]*kernel[1]+tmp[8698]*kernel[2]+tmp[8796]*kernel[3]+tmp[8797]*kernel[4]+tmp[8798]*kernel[5]+tmp[8896]*kernel[6]+tmp[8897]*kernel[7]+tmp[8898]*kernel[8];
				ans[8798]<=tmp[8697]*kernel[0]+tmp[8698]*kernel[1]+tmp[8699]*kernel[2]+tmp[8797]*kernel[3]+tmp[8798]*kernel[4]+tmp[8799]*kernel[5]+tmp[8897]*kernel[6]+tmp[8898]*kernel[7]+tmp[8899]*kernel[8];
				ans[8799]<=tmp[8698]*kernel[0]+tmp[8699]*kernel[1]+tmp[8798]*kernel[3]+tmp[8799]*kernel[4]+tmp[8898]*kernel[6]+tmp[8899]*kernel[7];
				ans[8800]<=tmp[8700]*kernel[1]+tmp[8701]*kernel[2]+tmp[8800]*kernel[4]+tmp[8801]*kernel[5]+tmp[8900]*kernel[7]+tmp[8901]*kernel[8];
				ans[8801]<=tmp[8700]*kernel[0]+tmp[8701]*kernel[1]+tmp[8702]*kernel[2]+tmp[8800]*kernel[3]+tmp[8801]*kernel[4]+tmp[8802]*kernel[5]+tmp[8900]*kernel[6]+tmp[8901]*kernel[7]+tmp[8902]*kernel[8];
				ans[8802]<=tmp[8701]*kernel[0]+tmp[8702]*kernel[1]+tmp[8703]*kernel[2]+tmp[8801]*kernel[3]+tmp[8802]*kernel[4]+tmp[8803]*kernel[5]+tmp[8901]*kernel[6]+tmp[8902]*kernel[7]+tmp[8903]*kernel[8];
				ans[8803]<=tmp[8702]*kernel[0]+tmp[8703]*kernel[1]+tmp[8704]*kernel[2]+tmp[8802]*kernel[3]+tmp[8803]*kernel[4]+tmp[8804]*kernel[5]+tmp[8902]*kernel[6]+tmp[8903]*kernel[7]+tmp[8904]*kernel[8];
				ans[8804]<=tmp[8703]*kernel[0]+tmp[8704]*kernel[1]+tmp[8705]*kernel[2]+tmp[8803]*kernel[3]+tmp[8804]*kernel[4]+tmp[8805]*kernel[5]+tmp[8903]*kernel[6]+tmp[8904]*kernel[7]+tmp[8905]*kernel[8];
				ans[8805]<=tmp[8704]*kernel[0]+tmp[8705]*kernel[1]+tmp[8706]*kernel[2]+tmp[8804]*kernel[3]+tmp[8805]*kernel[4]+tmp[8806]*kernel[5]+tmp[8904]*kernel[6]+tmp[8905]*kernel[7]+tmp[8906]*kernel[8];
				ans[8806]<=tmp[8705]*kernel[0]+tmp[8706]*kernel[1]+tmp[8707]*kernel[2]+tmp[8805]*kernel[3]+tmp[8806]*kernel[4]+tmp[8807]*kernel[5]+tmp[8905]*kernel[6]+tmp[8906]*kernel[7]+tmp[8907]*kernel[8];
				ans[8807]<=tmp[8706]*kernel[0]+tmp[8707]*kernel[1]+tmp[8708]*kernel[2]+tmp[8806]*kernel[3]+tmp[8807]*kernel[4]+tmp[8808]*kernel[5]+tmp[8906]*kernel[6]+tmp[8907]*kernel[7]+tmp[8908]*kernel[8];
				ans[8808]<=tmp[8707]*kernel[0]+tmp[8708]*kernel[1]+tmp[8709]*kernel[2]+tmp[8807]*kernel[3]+tmp[8808]*kernel[4]+tmp[8809]*kernel[5]+tmp[8907]*kernel[6]+tmp[8908]*kernel[7]+tmp[8909]*kernel[8];
				ans[8809]<=tmp[8708]*kernel[0]+tmp[8709]*kernel[1]+tmp[8710]*kernel[2]+tmp[8808]*kernel[3]+tmp[8809]*kernel[4]+tmp[8810]*kernel[5]+tmp[8908]*kernel[6]+tmp[8909]*kernel[7]+tmp[8910]*kernel[8];
				ans[8810]<=tmp[8709]*kernel[0]+tmp[8710]*kernel[1]+tmp[8711]*kernel[2]+tmp[8809]*kernel[3]+tmp[8810]*kernel[4]+tmp[8811]*kernel[5]+tmp[8909]*kernel[6]+tmp[8910]*kernel[7]+tmp[8911]*kernel[8];
				ans[8811]<=tmp[8710]*kernel[0]+tmp[8711]*kernel[1]+tmp[8712]*kernel[2]+tmp[8810]*kernel[3]+tmp[8811]*kernel[4]+tmp[8812]*kernel[5]+tmp[8910]*kernel[6]+tmp[8911]*kernel[7]+tmp[8912]*kernel[8];
				ans[8812]<=tmp[8711]*kernel[0]+tmp[8712]*kernel[1]+tmp[8713]*kernel[2]+tmp[8811]*kernel[3]+tmp[8812]*kernel[4]+tmp[8813]*kernel[5]+tmp[8911]*kernel[6]+tmp[8912]*kernel[7]+tmp[8913]*kernel[8];
				ans[8813]<=tmp[8712]*kernel[0]+tmp[8713]*kernel[1]+tmp[8714]*kernel[2]+tmp[8812]*kernel[3]+tmp[8813]*kernel[4]+tmp[8814]*kernel[5]+tmp[8912]*kernel[6]+tmp[8913]*kernel[7]+tmp[8914]*kernel[8];
				ans[8814]<=tmp[8713]*kernel[0]+tmp[8714]*kernel[1]+tmp[8715]*kernel[2]+tmp[8813]*kernel[3]+tmp[8814]*kernel[4]+tmp[8815]*kernel[5]+tmp[8913]*kernel[6]+tmp[8914]*kernel[7]+tmp[8915]*kernel[8];
				ans[8815]<=tmp[8714]*kernel[0]+tmp[8715]*kernel[1]+tmp[8716]*kernel[2]+tmp[8814]*kernel[3]+tmp[8815]*kernel[4]+tmp[8816]*kernel[5]+tmp[8914]*kernel[6]+tmp[8915]*kernel[7]+tmp[8916]*kernel[8];
				ans[8816]<=tmp[8715]*kernel[0]+tmp[8716]*kernel[1]+tmp[8717]*kernel[2]+tmp[8815]*kernel[3]+tmp[8816]*kernel[4]+tmp[8817]*kernel[5]+tmp[8915]*kernel[6]+tmp[8916]*kernel[7]+tmp[8917]*kernel[8];
				ans[8817]<=tmp[8716]*kernel[0]+tmp[8717]*kernel[1]+tmp[8718]*kernel[2]+tmp[8816]*kernel[3]+tmp[8817]*kernel[4]+tmp[8818]*kernel[5]+tmp[8916]*kernel[6]+tmp[8917]*kernel[7]+tmp[8918]*kernel[8];
				ans[8818]<=tmp[8717]*kernel[0]+tmp[8718]*kernel[1]+tmp[8719]*kernel[2]+tmp[8817]*kernel[3]+tmp[8818]*kernel[4]+tmp[8819]*kernel[5]+tmp[8917]*kernel[6]+tmp[8918]*kernel[7]+tmp[8919]*kernel[8];
				ans[8819]<=tmp[8718]*kernel[0]+tmp[8719]*kernel[1]+tmp[8720]*kernel[2]+tmp[8818]*kernel[3]+tmp[8819]*kernel[4]+tmp[8820]*kernel[5]+tmp[8918]*kernel[6]+tmp[8919]*kernel[7]+tmp[8920]*kernel[8];
				ans[8820]<=tmp[8719]*kernel[0]+tmp[8720]*kernel[1]+tmp[8721]*kernel[2]+tmp[8819]*kernel[3]+tmp[8820]*kernel[4]+tmp[8821]*kernel[5]+tmp[8919]*kernel[6]+tmp[8920]*kernel[7]+tmp[8921]*kernel[8];
				ans[8821]<=tmp[8720]*kernel[0]+tmp[8721]*kernel[1]+tmp[8722]*kernel[2]+tmp[8820]*kernel[3]+tmp[8821]*kernel[4]+tmp[8822]*kernel[5]+tmp[8920]*kernel[6]+tmp[8921]*kernel[7]+tmp[8922]*kernel[8];
				ans[8822]<=tmp[8721]*kernel[0]+tmp[8722]*kernel[1]+tmp[8723]*kernel[2]+tmp[8821]*kernel[3]+tmp[8822]*kernel[4]+tmp[8823]*kernel[5]+tmp[8921]*kernel[6]+tmp[8922]*kernel[7]+tmp[8923]*kernel[8];
				ans[8823]<=tmp[8722]*kernel[0]+tmp[8723]*kernel[1]+tmp[8724]*kernel[2]+tmp[8822]*kernel[3]+tmp[8823]*kernel[4]+tmp[8824]*kernel[5]+tmp[8922]*kernel[6]+tmp[8923]*kernel[7]+tmp[8924]*kernel[8];
				ans[8824]<=tmp[8723]*kernel[0]+tmp[8724]*kernel[1]+tmp[8725]*kernel[2]+tmp[8823]*kernel[3]+tmp[8824]*kernel[4]+tmp[8825]*kernel[5]+tmp[8923]*kernel[6]+tmp[8924]*kernel[7]+tmp[8925]*kernel[8];
				ans[8825]<=tmp[8724]*kernel[0]+tmp[8725]*kernel[1]+tmp[8726]*kernel[2]+tmp[8824]*kernel[3]+tmp[8825]*kernel[4]+tmp[8826]*kernel[5]+tmp[8924]*kernel[6]+tmp[8925]*kernel[7]+tmp[8926]*kernel[8];
				ans[8826]<=tmp[8725]*kernel[0]+tmp[8726]*kernel[1]+tmp[8727]*kernel[2]+tmp[8825]*kernel[3]+tmp[8826]*kernel[4]+tmp[8827]*kernel[5]+tmp[8925]*kernel[6]+tmp[8926]*kernel[7]+tmp[8927]*kernel[8];
				ans[8827]<=tmp[8726]*kernel[0]+tmp[8727]*kernel[1]+tmp[8728]*kernel[2]+tmp[8826]*kernel[3]+tmp[8827]*kernel[4]+tmp[8828]*kernel[5]+tmp[8926]*kernel[6]+tmp[8927]*kernel[7]+tmp[8928]*kernel[8];
				ans[8828]<=tmp[8727]*kernel[0]+tmp[8728]*kernel[1]+tmp[8729]*kernel[2]+tmp[8827]*kernel[3]+tmp[8828]*kernel[4]+tmp[8829]*kernel[5]+tmp[8927]*kernel[6]+tmp[8928]*kernel[7]+tmp[8929]*kernel[8];
				ans[8829]<=tmp[8728]*kernel[0]+tmp[8729]*kernel[1]+tmp[8730]*kernel[2]+tmp[8828]*kernel[3]+tmp[8829]*kernel[4]+tmp[8830]*kernel[5]+tmp[8928]*kernel[6]+tmp[8929]*kernel[7]+tmp[8930]*kernel[8];
				ans[8830]<=tmp[8729]*kernel[0]+tmp[8730]*kernel[1]+tmp[8731]*kernel[2]+tmp[8829]*kernel[3]+tmp[8830]*kernel[4]+tmp[8831]*kernel[5]+tmp[8929]*kernel[6]+tmp[8930]*kernel[7]+tmp[8931]*kernel[8];
				ans[8831]<=tmp[8730]*kernel[0]+tmp[8731]*kernel[1]+tmp[8732]*kernel[2]+tmp[8830]*kernel[3]+tmp[8831]*kernel[4]+tmp[8832]*kernel[5]+tmp[8930]*kernel[6]+tmp[8931]*kernel[7]+tmp[8932]*kernel[8];
				ans[8832]<=tmp[8731]*kernel[0]+tmp[8732]*kernel[1]+tmp[8733]*kernel[2]+tmp[8831]*kernel[3]+tmp[8832]*kernel[4]+tmp[8833]*kernel[5]+tmp[8931]*kernel[6]+tmp[8932]*kernel[7]+tmp[8933]*kernel[8];
				ans[8833]<=tmp[8732]*kernel[0]+tmp[8733]*kernel[1]+tmp[8734]*kernel[2]+tmp[8832]*kernel[3]+tmp[8833]*kernel[4]+tmp[8834]*kernel[5]+tmp[8932]*kernel[6]+tmp[8933]*kernel[7]+tmp[8934]*kernel[8];
				ans[8834]<=tmp[8733]*kernel[0]+tmp[8734]*kernel[1]+tmp[8735]*kernel[2]+tmp[8833]*kernel[3]+tmp[8834]*kernel[4]+tmp[8835]*kernel[5]+tmp[8933]*kernel[6]+tmp[8934]*kernel[7]+tmp[8935]*kernel[8];
				ans[8835]<=tmp[8734]*kernel[0]+tmp[8735]*kernel[1]+tmp[8736]*kernel[2]+tmp[8834]*kernel[3]+tmp[8835]*kernel[4]+tmp[8836]*kernel[5]+tmp[8934]*kernel[6]+tmp[8935]*kernel[7]+tmp[8936]*kernel[8];
				ans[8836]<=tmp[8735]*kernel[0]+tmp[8736]*kernel[1]+tmp[8737]*kernel[2]+tmp[8835]*kernel[3]+tmp[8836]*kernel[4]+tmp[8837]*kernel[5]+tmp[8935]*kernel[6]+tmp[8936]*kernel[7]+tmp[8937]*kernel[8];
				ans[8837]<=tmp[8736]*kernel[0]+tmp[8737]*kernel[1]+tmp[8738]*kernel[2]+tmp[8836]*kernel[3]+tmp[8837]*kernel[4]+tmp[8838]*kernel[5]+tmp[8936]*kernel[6]+tmp[8937]*kernel[7]+tmp[8938]*kernel[8];
				ans[8838]<=tmp[8737]*kernel[0]+tmp[8738]*kernel[1]+tmp[8739]*kernel[2]+tmp[8837]*kernel[3]+tmp[8838]*kernel[4]+tmp[8839]*kernel[5]+tmp[8937]*kernel[6]+tmp[8938]*kernel[7]+tmp[8939]*kernel[8];
				ans[8839]<=tmp[8738]*kernel[0]+tmp[8739]*kernel[1]+tmp[8740]*kernel[2]+tmp[8838]*kernel[3]+tmp[8839]*kernel[4]+tmp[8840]*kernel[5]+tmp[8938]*kernel[6]+tmp[8939]*kernel[7]+tmp[8940]*kernel[8];
				ans[8840]<=tmp[8739]*kernel[0]+tmp[8740]*kernel[1]+tmp[8741]*kernel[2]+tmp[8839]*kernel[3]+tmp[8840]*kernel[4]+tmp[8841]*kernel[5]+tmp[8939]*kernel[6]+tmp[8940]*kernel[7]+tmp[8941]*kernel[8];
				ans[8841]<=tmp[8740]*kernel[0]+tmp[8741]*kernel[1]+tmp[8742]*kernel[2]+tmp[8840]*kernel[3]+tmp[8841]*kernel[4]+tmp[8842]*kernel[5]+tmp[8940]*kernel[6]+tmp[8941]*kernel[7]+tmp[8942]*kernel[8];
				ans[8842]<=tmp[8741]*kernel[0]+tmp[8742]*kernel[1]+tmp[8743]*kernel[2]+tmp[8841]*kernel[3]+tmp[8842]*kernel[4]+tmp[8843]*kernel[5]+tmp[8941]*kernel[6]+tmp[8942]*kernel[7]+tmp[8943]*kernel[8];
				ans[8843]<=tmp[8742]*kernel[0]+tmp[8743]*kernel[1]+tmp[8744]*kernel[2]+tmp[8842]*kernel[3]+tmp[8843]*kernel[4]+tmp[8844]*kernel[5]+tmp[8942]*kernel[6]+tmp[8943]*kernel[7]+tmp[8944]*kernel[8];
				ans[8844]<=tmp[8743]*kernel[0]+tmp[8744]*kernel[1]+tmp[8745]*kernel[2]+tmp[8843]*kernel[3]+tmp[8844]*kernel[4]+tmp[8845]*kernel[5]+tmp[8943]*kernel[6]+tmp[8944]*kernel[7]+tmp[8945]*kernel[8];
				ans[8845]<=tmp[8744]*kernel[0]+tmp[8745]*kernel[1]+tmp[8746]*kernel[2]+tmp[8844]*kernel[3]+tmp[8845]*kernel[4]+tmp[8846]*kernel[5]+tmp[8944]*kernel[6]+tmp[8945]*kernel[7]+tmp[8946]*kernel[8];
				ans[8846]<=tmp[8745]*kernel[0]+tmp[8746]*kernel[1]+tmp[8747]*kernel[2]+tmp[8845]*kernel[3]+tmp[8846]*kernel[4]+tmp[8847]*kernel[5]+tmp[8945]*kernel[6]+tmp[8946]*kernel[7]+tmp[8947]*kernel[8];
				ans[8847]<=tmp[8746]*kernel[0]+tmp[8747]*kernel[1]+tmp[8748]*kernel[2]+tmp[8846]*kernel[3]+tmp[8847]*kernel[4]+tmp[8848]*kernel[5]+tmp[8946]*kernel[6]+tmp[8947]*kernel[7]+tmp[8948]*kernel[8];
				ans[8848]<=tmp[8747]*kernel[0]+tmp[8748]*kernel[1]+tmp[8749]*kernel[2]+tmp[8847]*kernel[3]+tmp[8848]*kernel[4]+tmp[8849]*kernel[5]+tmp[8947]*kernel[6]+tmp[8948]*kernel[7]+tmp[8949]*kernel[8];
				ans[8849]<=tmp[8748]*kernel[0]+tmp[8749]*kernel[1]+tmp[8750]*kernel[2]+tmp[8848]*kernel[3]+tmp[8849]*kernel[4]+tmp[8850]*kernel[5]+tmp[8948]*kernel[6]+tmp[8949]*kernel[7]+tmp[8950]*kernel[8];
				ans[8850]<=tmp[8749]*kernel[0]+tmp[8750]*kernel[1]+tmp[8751]*kernel[2]+tmp[8849]*kernel[3]+tmp[8850]*kernel[4]+tmp[8851]*kernel[5]+tmp[8949]*kernel[6]+tmp[8950]*kernel[7]+tmp[8951]*kernel[8];
				ans[8851]<=tmp[8750]*kernel[0]+tmp[8751]*kernel[1]+tmp[8752]*kernel[2]+tmp[8850]*kernel[3]+tmp[8851]*kernel[4]+tmp[8852]*kernel[5]+tmp[8950]*kernel[6]+tmp[8951]*kernel[7]+tmp[8952]*kernel[8];
				ans[8852]<=tmp[8751]*kernel[0]+tmp[8752]*kernel[1]+tmp[8753]*kernel[2]+tmp[8851]*kernel[3]+tmp[8852]*kernel[4]+tmp[8853]*kernel[5]+tmp[8951]*kernel[6]+tmp[8952]*kernel[7]+tmp[8953]*kernel[8];
				ans[8853]<=tmp[8752]*kernel[0]+tmp[8753]*kernel[1]+tmp[8754]*kernel[2]+tmp[8852]*kernel[3]+tmp[8853]*kernel[4]+tmp[8854]*kernel[5]+tmp[8952]*kernel[6]+tmp[8953]*kernel[7]+tmp[8954]*kernel[8];
				ans[8854]<=tmp[8753]*kernel[0]+tmp[8754]*kernel[1]+tmp[8755]*kernel[2]+tmp[8853]*kernel[3]+tmp[8854]*kernel[4]+tmp[8855]*kernel[5]+tmp[8953]*kernel[6]+tmp[8954]*kernel[7]+tmp[8955]*kernel[8];
				ans[8855]<=tmp[8754]*kernel[0]+tmp[8755]*kernel[1]+tmp[8756]*kernel[2]+tmp[8854]*kernel[3]+tmp[8855]*kernel[4]+tmp[8856]*kernel[5]+tmp[8954]*kernel[6]+tmp[8955]*kernel[7]+tmp[8956]*kernel[8];
				ans[8856]<=tmp[8755]*kernel[0]+tmp[8756]*kernel[1]+tmp[8757]*kernel[2]+tmp[8855]*kernel[3]+tmp[8856]*kernel[4]+tmp[8857]*kernel[5]+tmp[8955]*kernel[6]+tmp[8956]*kernel[7]+tmp[8957]*kernel[8];
				ans[8857]<=tmp[8756]*kernel[0]+tmp[8757]*kernel[1]+tmp[8758]*kernel[2]+tmp[8856]*kernel[3]+tmp[8857]*kernel[4]+tmp[8858]*kernel[5]+tmp[8956]*kernel[6]+tmp[8957]*kernel[7]+tmp[8958]*kernel[8];
				ans[8858]<=tmp[8757]*kernel[0]+tmp[8758]*kernel[1]+tmp[8759]*kernel[2]+tmp[8857]*kernel[3]+tmp[8858]*kernel[4]+tmp[8859]*kernel[5]+tmp[8957]*kernel[6]+tmp[8958]*kernel[7]+tmp[8959]*kernel[8];
				ans[8859]<=tmp[8758]*kernel[0]+tmp[8759]*kernel[1]+tmp[8760]*kernel[2]+tmp[8858]*kernel[3]+tmp[8859]*kernel[4]+tmp[8860]*kernel[5]+tmp[8958]*kernel[6]+tmp[8959]*kernel[7]+tmp[8960]*kernel[8];
				ans[8860]<=tmp[8759]*kernel[0]+tmp[8760]*kernel[1]+tmp[8761]*kernel[2]+tmp[8859]*kernel[3]+tmp[8860]*kernel[4]+tmp[8861]*kernel[5]+tmp[8959]*kernel[6]+tmp[8960]*kernel[7]+tmp[8961]*kernel[8];
				ans[8861]<=tmp[8760]*kernel[0]+tmp[8761]*kernel[1]+tmp[8762]*kernel[2]+tmp[8860]*kernel[3]+tmp[8861]*kernel[4]+tmp[8862]*kernel[5]+tmp[8960]*kernel[6]+tmp[8961]*kernel[7]+tmp[8962]*kernel[8];
				ans[8862]<=tmp[8761]*kernel[0]+tmp[8762]*kernel[1]+tmp[8763]*kernel[2]+tmp[8861]*kernel[3]+tmp[8862]*kernel[4]+tmp[8863]*kernel[5]+tmp[8961]*kernel[6]+tmp[8962]*kernel[7]+tmp[8963]*kernel[8];
				ans[8863]<=tmp[8762]*kernel[0]+tmp[8763]*kernel[1]+tmp[8764]*kernel[2]+tmp[8862]*kernel[3]+tmp[8863]*kernel[4]+tmp[8864]*kernel[5]+tmp[8962]*kernel[6]+tmp[8963]*kernel[7]+tmp[8964]*kernel[8];
				ans[8864]<=tmp[8763]*kernel[0]+tmp[8764]*kernel[1]+tmp[8765]*kernel[2]+tmp[8863]*kernel[3]+tmp[8864]*kernel[4]+tmp[8865]*kernel[5]+tmp[8963]*kernel[6]+tmp[8964]*kernel[7]+tmp[8965]*kernel[8];
				ans[8865]<=tmp[8764]*kernel[0]+tmp[8765]*kernel[1]+tmp[8766]*kernel[2]+tmp[8864]*kernel[3]+tmp[8865]*kernel[4]+tmp[8866]*kernel[5]+tmp[8964]*kernel[6]+tmp[8965]*kernel[7]+tmp[8966]*kernel[8];
				ans[8866]<=tmp[8765]*kernel[0]+tmp[8766]*kernel[1]+tmp[8767]*kernel[2]+tmp[8865]*kernel[3]+tmp[8866]*kernel[4]+tmp[8867]*kernel[5]+tmp[8965]*kernel[6]+tmp[8966]*kernel[7]+tmp[8967]*kernel[8];
				ans[8867]<=tmp[8766]*kernel[0]+tmp[8767]*kernel[1]+tmp[8768]*kernel[2]+tmp[8866]*kernel[3]+tmp[8867]*kernel[4]+tmp[8868]*kernel[5]+tmp[8966]*kernel[6]+tmp[8967]*kernel[7]+tmp[8968]*kernel[8];
				ans[8868]<=tmp[8767]*kernel[0]+tmp[8768]*kernel[1]+tmp[8769]*kernel[2]+tmp[8867]*kernel[3]+tmp[8868]*kernel[4]+tmp[8869]*kernel[5]+tmp[8967]*kernel[6]+tmp[8968]*kernel[7]+tmp[8969]*kernel[8];
				ans[8869]<=tmp[8768]*kernel[0]+tmp[8769]*kernel[1]+tmp[8770]*kernel[2]+tmp[8868]*kernel[3]+tmp[8869]*kernel[4]+tmp[8870]*kernel[5]+tmp[8968]*kernel[6]+tmp[8969]*kernel[7]+tmp[8970]*kernel[8];
				ans[8870]<=tmp[8769]*kernel[0]+tmp[8770]*kernel[1]+tmp[8771]*kernel[2]+tmp[8869]*kernel[3]+tmp[8870]*kernel[4]+tmp[8871]*kernel[5]+tmp[8969]*kernel[6]+tmp[8970]*kernel[7]+tmp[8971]*kernel[8];
				ans[8871]<=tmp[8770]*kernel[0]+tmp[8771]*kernel[1]+tmp[8772]*kernel[2]+tmp[8870]*kernel[3]+tmp[8871]*kernel[4]+tmp[8872]*kernel[5]+tmp[8970]*kernel[6]+tmp[8971]*kernel[7]+tmp[8972]*kernel[8];
				ans[8872]<=tmp[8771]*kernel[0]+tmp[8772]*kernel[1]+tmp[8773]*kernel[2]+tmp[8871]*kernel[3]+tmp[8872]*kernel[4]+tmp[8873]*kernel[5]+tmp[8971]*kernel[6]+tmp[8972]*kernel[7]+tmp[8973]*kernel[8];
				ans[8873]<=tmp[8772]*kernel[0]+tmp[8773]*kernel[1]+tmp[8774]*kernel[2]+tmp[8872]*kernel[3]+tmp[8873]*kernel[4]+tmp[8874]*kernel[5]+tmp[8972]*kernel[6]+tmp[8973]*kernel[7]+tmp[8974]*kernel[8];
				ans[8874]<=tmp[8773]*kernel[0]+tmp[8774]*kernel[1]+tmp[8775]*kernel[2]+tmp[8873]*kernel[3]+tmp[8874]*kernel[4]+tmp[8875]*kernel[5]+tmp[8973]*kernel[6]+tmp[8974]*kernel[7]+tmp[8975]*kernel[8];
				ans[8875]<=tmp[8774]*kernel[0]+tmp[8775]*kernel[1]+tmp[8776]*kernel[2]+tmp[8874]*kernel[3]+tmp[8875]*kernel[4]+tmp[8876]*kernel[5]+tmp[8974]*kernel[6]+tmp[8975]*kernel[7]+tmp[8976]*kernel[8];
				ans[8876]<=tmp[8775]*kernel[0]+tmp[8776]*kernel[1]+tmp[8777]*kernel[2]+tmp[8875]*kernel[3]+tmp[8876]*kernel[4]+tmp[8877]*kernel[5]+tmp[8975]*kernel[6]+tmp[8976]*kernel[7]+tmp[8977]*kernel[8];
				ans[8877]<=tmp[8776]*kernel[0]+tmp[8777]*kernel[1]+tmp[8778]*kernel[2]+tmp[8876]*kernel[3]+tmp[8877]*kernel[4]+tmp[8878]*kernel[5]+tmp[8976]*kernel[6]+tmp[8977]*kernel[7]+tmp[8978]*kernel[8];
				ans[8878]<=tmp[8777]*kernel[0]+tmp[8778]*kernel[1]+tmp[8779]*kernel[2]+tmp[8877]*kernel[3]+tmp[8878]*kernel[4]+tmp[8879]*kernel[5]+tmp[8977]*kernel[6]+tmp[8978]*kernel[7]+tmp[8979]*kernel[8];
				ans[8879]<=tmp[8778]*kernel[0]+tmp[8779]*kernel[1]+tmp[8780]*kernel[2]+tmp[8878]*kernel[3]+tmp[8879]*kernel[4]+tmp[8880]*kernel[5]+tmp[8978]*kernel[6]+tmp[8979]*kernel[7]+tmp[8980]*kernel[8];
				ans[8880]<=tmp[8779]*kernel[0]+tmp[8780]*kernel[1]+tmp[8781]*kernel[2]+tmp[8879]*kernel[3]+tmp[8880]*kernel[4]+tmp[8881]*kernel[5]+tmp[8979]*kernel[6]+tmp[8980]*kernel[7]+tmp[8981]*kernel[8];
				ans[8881]<=tmp[8780]*kernel[0]+tmp[8781]*kernel[1]+tmp[8782]*kernel[2]+tmp[8880]*kernel[3]+tmp[8881]*kernel[4]+tmp[8882]*kernel[5]+tmp[8980]*kernel[6]+tmp[8981]*kernel[7]+tmp[8982]*kernel[8];
				ans[8882]<=tmp[8781]*kernel[0]+tmp[8782]*kernel[1]+tmp[8783]*kernel[2]+tmp[8881]*kernel[3]+tmp[8882]*kernel[4]+tmp[8883]*kernel[5]+tmp[8981]*kernel[6]+tmp[8982]*kernel[7]+tmp[8983]*kernel[8];
				ans[8883]<=tmp[8782]*kernel[0]+tmp[8783]*kernel[1]+tmp[8784]*kernel[2]+tmp[8882]*kernel[3]+tmp[8883]*kernel[4]+tmp[8884]*kernel[5]+tmp[8982]*kernel[6]+tmp[8983]*kernel[7]+tmp[8984]*kernel[8];
				ans[8884]<=tmp[8783]*kernel[0]+tmp[8784]*kernel[1]+tmp[8785]*kernel[2]+tmp[8883]*kernel[3]+tmp[8884]*kernel[4]+tmp[8885]*kernel[5]+tmp[8983]*kernel[6]+tmp[8984]*kernel[7]+tmp[8985]*kernel[8];
				ans[8885]<=tmp[8784]*kernel[0]+tmp[8785]*kernel[1]+tmp[8786]*kernel[2]+tmp[8884]*kernel[3]+tmp[8885]*kernel[4]+tmp[8886]*kernel[5]+tmp[8984]*kernel[6]+tmp[8985]*kernel[7]+tmp[8986]*kernel[8];
				ans[8886]<=tmp[8785]*kernel[0]+tmp[8786]*kernel[1]+tmp[8787]*kernel[2]+tmp[8885]*kernel[3]+tmp[8886]*kernel[4]+tmp[8887]*kernel[5]+tmp[8985]*kernel[6]+tmp[8986]*kernel[7]+tmp[8987]*kernel[8];
				ans[8887]<=tmp[8786]*kernel[0]+tmp[8787]*kernel[1]+tmp[8788]*kernel[2]+tmp[8886]*kernel[3]+tmp[8887]*kernel[4]+tmp[8888]*kernel[5]+tmp[8986]*kernel[6]+tmp[8987]*kernel[7]+tmp[8988]*kernel[8];
				ans[8888]<=tmp[8787]*kernel[0]+tmp[8788]*kernel[1]+tmp[8789]*kernel[2]+tmp[8887]*kernel[3]+tmp[8888]*kernel[4]+tmp[8889]*kernel[5]+tmp[8987]*kernel[6]+tmp[8988]*kernel[7]+tmp[8989]*kernel[8];
				ans[8889]<=tmp[8788]*kernel[0]+tmp[8789]*kernel[1]+tmp[8790]*kernel[2]+tmp[8888]*kernel[3]+tmp[8889]*kernel[4]+tmp[8890]*kernel[5]+tmp[8988]*kernel[6]+tmp[8989]*kernel[7]+tmp[8990]*kernel[8];
				ans[8890]<=tmp[8789]*kernel[0]+tmp[8790]*kernel[1]+tmp[8791]*kernel[2]+tmp[8889]*kernel[3]+tmp[8890]*kernel[4]+tmp[8891]*kernel[5]+tmp[8989]*kernel[6]+tmp[8990]*kernel[7]+tmp[8991]*kernel[8];
				ans[8891]<=tmp[8790]*kernel[0]+tmp[8791]*kernel[1]+tmp[8792]*kernel[2]+tmp[8890]*kernel[3]+tmp[8891]*kernel[4]+tmp[8892]*kernel[5]+tmp[8990]*kernel[6]+tmp[8991]*kernel[7]+tmp[8992]*kernel[8];
				ans[8892]<=tmp[8791]*kernel[0]+tmp[8792]*kernel[1]+tmp[8793]*kernel[2]+tmp[8891]*kernel[3]+tmp[8892]*kernel[4]+tmp[8893]*kernel[5]+tmp[8991]*kernel[6]+tmp[8992]*kernel[7]+tmp[8993]*kernel[8];
				ans[8893]<=tmp[8792]*kernel[0]+tmp[8793]*kernel[1]+tmp[8794]*kernel[2]+tmp[8892]*kernel[3]+tmp[8893]*kernel[4]+tmp[8894]*kernel[5]+tmp[8992]*kernel[6]+tmp[8993]*kernel[7]+tmp[8994]*kernel[8];
				ans[8894]<=tmp[8793]*kernel[0]+tmp[8794]*kernel[1]+tmp[8795]*kernel[2]+tmp[8893]*kernel[3]+tmp[8894]*kernel[4]+tmp[8895]*kernel[5]+tmp[8993]*kernel[6]+tmp[8994]*kernel[7]+tmp[8995]*kernel[8];
				ans[8895]<=tmp[8794]*kernel[0]+tmp[8795]*kernel[1]+tmp[8796]*kernel[2]+tmp[8894]*kernel[3]+tmp[8895]*kernel[4]+tmp[8896]*kernel[5]+tmp[8994]*kernel[6]+tmp[8995]*kernel[7]+tmp[8996]*kernel[8];
				ans[8896]<=tmp[8795]*kernel[0]+tmp[8796]*kernel[1]+tmp[8797]*kernel[2]+tmp[8895]*kernel[3]+tmp[8896]*kernel[4]+tmp[8897]*kernel[5]+tmp[8995]*kernel[6]+tmp[8996]*kernel[7]+tmp[8997]*kernel[8];
				ans[8897]<=tmp[8796]*kernel[0]+tmp[8797]*kernel[1]+tmp[8798]*kernel[2]+tmp[8896]*kernel[3]+tmp[8897]*kernel[4]+tmp[8898]*kernel[5]+tmp[8996]*kernel[6]+tmp[8997]*kernel[7]+tmp[8998]*kernel[8];
				ans[8898]<=tmp[8797]*kernel[0]+tmp[8798]*kernel[1]+tmp[8799]*kernel[2]+tmp[8897]*kernel[3]+tmp[8898]*kernel[4]+tmp[8899]*kernel[5]+tmp[8997]*kernel[6]+tmp[8998]*kernel[7]+tmp[8999]*kernel[8];
				ans[8899]<=tmp[8798]*kernel[0]+tmp[8799]*kernel[1]+tmp[8898]*kernel[3]+tmp[8899]*kernel[4]+tmp[8998]*kernel[6]+tmp[8999]*kernel[7];
				ans[8900]<=tmp[8800]*kernel[1]+tmp[8801]*kernel[2]+tmp[8900]*kernel[4]+tmp[8901]*kernel[5]+tmp[9000]*kernel[7]+tmp[9001]*kernel[8];
				ans[8901]<=tmp[8800]*kernel[0]+tmp[8801]*kernel[1]+tmp[8802]*kernel[2]+tmp[8900]*kernel[3]+tmp[8901]*kernel[4]+tmp[8902]*kernel[5]+tmp[9000]*kernel[6]+tmp[9001]*kernel[7]+tmp[9002]*kernel[8];
				ans[8902]<=tmp[8801]*kernel[0]+tmp[8802]*kernel[1]+tmp[8803]*kernel[2]+tmp[8901]*kernel[3]+tmp[8902]*kernel[4]+tmp[8903]*kernel[5]+tmp[9001]*kernel[6]+tmp[9002]*kernel[7]+tmp[9003]*kernel[8];
				ans[8903]<=tmp[8802]*kernel[0]+tmp[8803]*kernel[1]+tmp[8804]*kernel[2]+tmp[8902]*kernel[3]+tmp[8903]*kernel[4]+tmp[8904]*kernel[5]+tmp[9002]*kernel[6]+tmp[9003]*kernel[7]+tmp[9004]*kernel[8];
				ans[8904]<=tmp[8803]*kernel[0]+tmp[8804]*kernel[1]+tmp[8805]*kernel[2]+tmp[8903]*kernel[3]+tmp[8904]*kernel[4]+tmp[8905]*kernel[5]+tmp[9003]*kernel[6]+tmp[9004]*kernel[7]+tmp[9005]*kernel[8];
				ans[8905]<=tmp[8804]*kernel[0]+tmp[8805]*kernel[1]+tmp[8806]*kernel[2]+tmp[8904]*kernel[3]+tmp[8905]*kernel[4]+tmp[8906]*kernel[5]+tmp[9004]*kernel[6]+tmp[9005]*kernel[7]+tmp[9006]*kernel[8];
				ans[8906]<=tmp[8805]*kernel[0]+tmp[8806]*kernel[1]+tmp[8807]*kernel[2]+tmp[8905]*kernel[3]+tmp[8906]*kernel[4]+tmp[8907]*kernel[5]+tmp[9005]*kernel[6]+tmp[9006]*kernel[7]+tmp[9007]*kernel[8];
				ans[8907]<=tmp[8806]*kernel[0]+tmp[8807]*kernel[1]+tmp[8808]*kernel[2]+tmp[8906]*kernel[3]+tmp[8907]*kernel[4]+tmp[8908]*kernel[5]+tmp[9006]*kernel[6]+tmp[9007]*kernel[7]+tmp[9008]*kernel[8];
				ans[8908]<=tmp[8807]*kernel[0]+tmp[8808]*kernel[1]+tmp[8809]*kernel[2]+tmp[8907]*kernel[3]+tmp[8908]*kernel[4]+tmp[8909]*kernel[5]+tmp[9007]*kernel[6]+tmp[9008]*kernel[7]+tmp[9009]*kernel[8];
				ans[8909]<=tmp[8808]*kernel[0]+tmp[8809]*kernel[1]+tmp[8810]*kernel[2]+tmp[8908]*kernel[3]+tmp[8909]*kernel[4]+tmp[8910]*kernel[5]+tmp[9008]*kernel[6]+tmp[9009]*kernel[7]+tmp[9010]*kernel[8];
				ans[8910]<=tmp[8809]*kernel[0]+tmp[8810]*kernel[1]+tmp[8811]*kernel[2]+tmp[8909]*kernel[3]+tmp[8910]*kernel[4]+tmp[8911]*kernel[5]+tmp[9009]*kernel[6]+tmp[9010]*kernel[7]+tmp[9011]*kernel[8];
				ans[8911]<=tmp[8810]*kernel[0]+tmp[8811]*kernel[1]+tmp[8812]*kernel[2]+tmp[8910]*kernel[3]+tmp[8911]*kernel[4]+tmp[8912]*kernel[5]+tmp[9010]*kernel[6]+tmp[9011]*kernel[7]+tmp[9012]*kernel[8];
				ans[8912]<=tmp[8811]*kernel[0]+tmp[8812]*kernel[1]+tmp[8813]*kernel[2]+tmp[8911]*kernel[3]+tmp[8912]*kernel[4]+tmp[8913]*kernel[5]+tmp[9011]*kernel[6]+tmp[9012]*kernel[7]+tmp[9013]*kernel[8];
				ans[8913]<=tmp[8812]*kernel[0]+tmp[8813]*kernel[1]+tmp[8814]*kernel[2]+tmp[8912]*kernel[3]+tmp[8913]*kernel[4]+tmp[8914]*kernel[5]+tmp[9012]*kernel[6]+tmp[9013]*kernel[7]+tmp[9014]*kernel[8];
				ans[8914]<=tmp[8813]*kernel[0]+tmp[8814]*kernel[1]+tmp[8815]*kernel[2]+tmp[8913]*kernel[3]+tmp[8914]*kernel[4]+tmp[8915]*kernel[5]+tmp[9013]*kernel[6]+tmp[9014]*kernel[7]+tmp[9015]*kernel[8];
				ans[8915]<=tmp[8814]*kernel[0]+tmp[8815]*kernel[1]+tmp[8816]*kernel[2]+tmp[8914]*kernel[3]+tmp[8915]*kernel[4]+tmp[8916]*kernel[5]+tmp[9014]*kernel[6]+tmp[9015]*kernel[7]+tmp[9016]*kernel[8];
				ans[8916]<=tmp[8815]*kernel[0]+tmp[8816]*kernel[1]+tmp[8817]*kernel[2]+tmp[8915]*kernel[3]+tmp[8916]*kernel[4]+tmp[8917]*kernel[5]+tmp[9015]*kernel[6]+tmp[9016]*kernel[7]+tmp[9017]*kernel[8];
				ans[8917]<=tmp[8816]*kernel[0]+tmp[8817]*kernel[1]+tmp[8818]*kernel[2]+tmp[8916]*kernel[3]+tmp[8917]*kernel[4]+tmp[8918]*kernel[5]+tmp[9016]*kernel[6]+tmp[9017]*kernel[7]+tmp[9018]*kernel[8];
				ans[8918]<=tmp[8817]*kernel[0]+tmp[8818]*kernel[1]+tmp[8819]*kernel[2]+tmp[8917]*kernel[3]+tmp[8918]*kernel[4]+tmp[8919]*kernel[5]+tmp[9017]*kernel[6]+tmp[9018]*kernel[7]+tmp[9019]*kernel[8];
				ans[8919]<=tmp[8818]*kernel[0]+tmp[8819]*kernel[1]+tmp[8820]*kernel[2]+tmp[8918]*kernel[3]+tmp[8919]*kernel[4]+tmp[8920]*kernel[5]+tmp[9018]*kernel[6]+tmp[9019]*kernel[7]+tmp[9020]*kernel[8];
				ans[8920]<=tmp[8819]*kernel[0]+tmp[8820]*kernel[1]+tmp[8821]*kernel[2]+tmp[8919]*kernel[3]+tmp[8920]*kernel[4]+tmp[8921]*kernel[5]+tmp[9019]*kernel[6]+tmp[9020]*kernel[7]+tmp[9021]*kernel[8];
				ans[8921]<=tmp[8820]*kernel[0]+tmp[8821]*kernel[1]+tmp[8822]*kernel[2]+tmp[8920]*kernel[3]+tmp[8921]*kernel[4]+tmp[8922]*kernel[5]+tmp[9020]*kernel[6]+tmp[9021]*kernel[7]+tmp[9022]*kernel[8];
				ans[8922]<=tmp[8821]*kernel[0]+tmp[8822]*kernel[1]+tmp[8823]*kernel[2]+tmp[8921]*kernel[3]+tmp[8922]*kernel[4]+tmp[8923]*kernel[5]+tmp[9021]*kernel[6]+tmp[9022]*kernel[7]+tmp[9023]*kernel[8];
				ans[8923]<=tmp[8822]*kernel[0]+tmp[8823]*kernel[1]+tmp[8824]*kernel[2]+tmp[8922]*kernel[3]+tmp[8923]*kernel[4]+tmp[8924]*kernel[5]+tmp[9022]*kernel[6]+tmp[9023]*kernel[7]+tmp[9024]*kernel[8];
				ans[8924]<=tmp[8823]*kernel[0]+tmp[8824]*kernel[1]+tmp[8825]*kernel[2]+tmp[8923]*kernel[3]+tmp[8924]*kernel[4]+tmp[8925]*kernel[5]+tmp[9023]*kernel[6]+tmp[9024]*kernel[7]+tmp[9025]*kernel[8];
				ans[8925]<=tmp[8824]*kernel[0]+tmp[8825]*kernel[1]+tmp[8826]*kernel[2]+tmp[8924]*kernel[3]+tmp[8925]*kernel[4]+tmp[8926]*kernel[5]+tmp[9024]*kernel[6]+tmp[9025]*kernel[7]+tmp[9026]*kernel[8];
				ans[8926]<=tmp[8825]*kernel[0]+tmp[8826]*kernel[1]+tmp[8827]*kernel[2]+tmp[8925]*kernel[3]+tmp[8926]*kernel[4]+tmp[8927]*kernel[5]+tmp[9025]*kernel[6]+tmp[9026]*kernel[7]+tmp[9027]*kernel[8];
				ans[8927]<=tmp[8826]*kernel[0]+tmp[8827]*kernel[1]+tmp[8828]*kernel[2]+tmp[8926]*kernel[3]+tmp[8927]*kernel[4]+tmp[8928]*kernel[5]+tmp[9026]*kernel[6]+tmp[9027]*kernel[7]+tmp[9028]*kernel[8];
				ans[8928]<=tmp[8827]*kernel[0]+tmp[8828]*kernel[1]+tmp[8829]*kernel[2]+tmp[8927]*kernel[3]+tmp[8928]*kernel[4]+tmp[8929]*kernel[5]+tmp[9027]*kernel[6]+tmp[9028]*kernel[7]+tmp[9029]*kernel[8];
				ans[8929]<=tmp[8828]*kernel[0]+tmp[8829]*kernel[1]+tmp[8830]*kernel[2]+tmp[8928]*kernel[3]+tmp[8929]*kernel[4]+tmp[8930]*kernel[5]+tmp[9028]*kernel[6]+tmp[9029]*kernel[7]+tmp[9030]*kernel[8];
				ans[8930]<=tmp[8829]*kernel[0]+tmp[8830]*kernel[1]+tmp[8831]*kernel[2]+tmp[8929]*kernel[3]+tmp[8930]*kernel[4]+tmp[8931]*kernel[5]+tmp[9029]*kernel[6]+tmp[9030]*kernel[7]+tmp[9031]*kernel[8];
				ans[8931]<=tmp[8830]*kernel[0]+tmp[8831]*kernel[1]+tmp[8832]*kernel[2]+tmp[8930]*kernel[3]+tmp[8931]*kernel[4]+tmp[8932]*kernel[5]+tmp[9030]*kernel[6]+tmp[9031]*kernel[7]+tmp[9032]*kernel[8];
				ans[8932]<=tmp[8831]*kernel[0]+tmp[8832]*kernel[1]+tmp[8833]*kernel[2]+tmp[8931]*kernel[3]+tmp[8932]*kernel[4]+tmp[8933]*kernel[5]+tmp[9031]*kernel[6]+tmp[9032]*kernel[7]+tmp[9033]*kernel[8];
				ans[8933]<=tmp[8832]*kernel[0]+tmp[8833]*kernel[1]+tmp[8834]*kernel[2]+tmp[8932]*kernel[3]+tmp[8933]*kernel[4]+tmp[8934]*kernel[5]+tmp[9032]*kernel[6]+tmp[9033]*kernel[7]+tmp[9034]*kernel[8];
				ans[8934]<=tmp[8833]*kernel[0]+tmp[8834]*kernel[1]+tmp[8835]*kernel[2]+tmp[8933]*kernel[3]+tmp[8934]*kernel[4]+tmp[8935]*kernel[5]+tmp[9033]*kernel[6]+tmp[9034]*kernel[7]+tmp[9035]*kernel[8];
				ans[8935]<=tmp[8834]*kernel[0]+tmp[8835]*kernel[1]+tmp[8836]*kernel[2]+tmp[8934]*kernel[3]+tmp[8935]*kernel[4]+tmp[8936]*kernel[5]+tmp[9034]*kernel[6]+tmp[9035]*kernel[7]+tmp[9036]*kernel[8];
				ans[8936]<=tmp[8835]*kernel[0]+tmp[8836]*kernel[1]+tmp[8837]*kernel[2]+tmp[8935]*kernel[3]+tmp[8936]*kernel[4]+tmp[8937]*kernel[5]+tmp[9035]*kernel[6]+tmp[9036]*kernel[7]+tmp[9037]*kernel[8];
				ans[8937]<=tmp[8836]*kernel[0]+tmp[8837]*kernel[1]+tmp[8838]*kernel[2]+tmp[8936]*kernel[3]+tmp[8937]*kernel[4]+tmp[8938]*kernel[5]+tmp[9036]*kernel[6]+tmp[9037]*kernel[7]+tmp[9038]*kernel[8];
				ans[8938]<=tmp[8837]*kernel[0]+tmp[8838]*kernel[1]+tmp[8839]*kernel[2]+tmp[8937]*kernel[3]+tmp[8938]*kernel[4]+tmp[8939]*kernel[5]+tmp[9037]*kernel[6]+tmp[9038]*kernel[7]+tmp[9039]*kernel[8];
				ans[8939]<=tmp[8838]*kernel[0]+tmp[8839]*kernel[1]+tmp[8840]*kernel[2]+tmp[8938]*kernel[3]+tmp[8939]*kernel[4]+tmp[8940]*kernel[5]+tmp[9038]*kernel[6]+tmp[9039]*kernel[7]+tmp[9040]*kernel[8];
				ans[8940]<=tmp[8839]*kernel[0]+tmp[8840]*kernel[1]+tmp[8841]*kernel[2]+tmp[8939]*kernel[3]+tmp[8940]*kernel[4]+tmp[8941]*kernel[5]+tmp[9039]*kernel[6]+tmp[9040]*kernel[7]+tmp[9041]*kernel[8];
				ans[8941]<=tmp[8840]*kernel[0]+tmp[8841]*kernel[1]+tmp[8842]*kernel[2]+tmp[8940]*kernel[3]+tmp[8941]*kernel[4]+tmp[8942]*kernel[5]+tmp[9040]*kernel[6]+tmp[9041]*kernel[7]+tmp[9042]*kernel[8];
				ans[8942]<=tmp[8841]*kernel[0]+tmp[8842]*kernel[1]+tmp[8843]*kernel[2]+tmp[8941]*kernel[3]+tmp[8942]*kernel[4]+tmp[8943]*kernel[5]+tmp[9041]*kernel[6]+tmp[9042]*kernel[7]+tmp[9043]*kernel[8];
				ans[8943]<=tmp[8842]*kernel[0]+tmp[8843]*kernel[1]+tmp[8844]*kernel[2]+tmp[8942]*kernel[3]+tmp[8943]*kernel[4]+tmp[8944]*kernel[5]+tmp[9042]*kernel[6]+tmp[9043]*kernel[7]+tmp[9044]*kernel[8];
				ans[8944]<=tmp[8843]*kernel[0]+tmp[8844]*kernel[1]+tmp[8845]*kernel[2]+tmp[8943]*kernel[3]+tmp[8944]*kernel[4]+tmp[8945]*kernel[5]+tmp[9043]*kernel[6]+tmp[9044]*kernel[7]+tmp[9045]*kernel[8];
				ans[8945]<=tmp[8844]*kernel[0]+tmp[8845]*kernel[1]+tmp[8846]*kernel[2]+tmp[8944]*kernel[3]+tmp[8945]*kernel[4]+tmp[8946]*kernel[5]+tmp[9044]*kernel[6]+tmp[9045]*kernel[7]+tmp[9046]*kernel[8];
				ans[8946]<=tmp[8845]*kernel[0]+tmp[8846]*kernel[1]+tmp[8847]*kernel[2]+tmp[8945]*kernel[3]+tmp[8946]*kernel[4]+tmp[8947]*kernel[5]+tmp[9045]*kernel[6]+tmp[9046]*kernel[7]+tmp[9047]*kernel[8];
				ans[8947]<=tmp[8846]*kernel[0]+tmp[8847]*kernel[1]+tmp[8848]*kernel[2]+tmp[8946]*kernel[3]+tmp[8947]*kernel[4]+tmp[8948]*kernel[5]+tmp[9046]*kernel[6]+tmp[9047]*kernel[7]+tmp[9048]*kernel[8];
				ans[8948]<=tmp[8847]*kernel[0]+tmp[8848]*kernel[1]+tmp[8849]*kernel[2]+tmp[8947]*kernel[3]+tmp[8948]*kernel[4]+tmp[8949]*kernel[5]+tmp[9047]*kernel[6]+tmp[9048]*kernel[7]+tmp[9049]*kernel[8];
				ans[8949]<=tmp[8848]*kernel[0]+tmp[8849]*kernel[1]+tmp[8850]*kernel[2]+tmp[8948]*kernel[3]+tmp[8949]*kernel[4]+tmp[8950]*kernel[5]+tmp[9048]*kernel[6]+tmp[9049]*kernel[7]+tmp[9050]*kernel[8];
				ans[8950]<=tmp[8849]*kernel[0]+tmp[8850]*kernel[1]+tmp[8851]*kernel[2]+tmp[8949]*kernel[3]+tmp[8950]*kernel[4]+tmp[8951]*kernel[5]+tmp[9049]*kernel[6]+tmp[9050]*kernel[7]+tmp[9051]*kernel[8];
				ans[8951]<=tmp[8850]*kernel[0]+tmp[8851]*kernel[1]+tmp[8852]*kernel[2]+tmp[8950]*kernel[3]+tmp[8951]*kernel[4]+tmp[8952]*kernel[5]+tmp[9050]*kernel[6]+tmp[9051]*kernel[7]+tmp[9052]*kernel[8];
				ans[8952]<=tmp[8851]*kernel[0]+tmp[8852]*kernel[1]+tmp[8853]*kernel[2]+tmp[8951]*kernel[3]+tmp[8952]*kernel[4]+tmp[8953]*kernel[5]+tmp[9051]*kernel[6]+tmp[9052]*kernel[7]+tmp[9053]*kernel[8];
				ans[8953]<=tmp[8852]*kernel[0]+tmp[8853]*kernel[1]+tmp[8854]*kernel[2]+tmp[8952]*kernel[3]+tmp[8953]*kernel[4]+tmp[8954]*kernel[5]+tmp[9052]*kernel[6]+tmp[9053]*kernel[7]+tmp[9054]*kernel[8];
				ans[8954]<=tmp[8853]*kernel[0]+tmp[8854]*kernel[1]+tmp[8855]*kernel[2]+tmp[8953]*kernel[3]+tmp[8954]*kernel[4]+tmp[8955]*kernel[5]+tmp[9053]*kernel[6]+tmp[9054]*kernel[7]+tmp[9055]*kernel[8];
				ans[8955]<=tmp[8854]*kernel[0]+tmp[8855]*kernel[1]+tmp[8856]*kernel[2]+tmp[8954]*kernel[3]+tmp[8955]*kernel[4]+tmp[8956]*kernel[5]+tmp[9054]*kernel[6]+tmp[9055]*kernel[7]+tmp[9056]*kernel[8];
				ans[8956]<=tmp[8855]*kernel[0]+tmp[8856]*kernel[1]+tmp[8857]*kernel[2]+tmp[8955]*kernel[3]+tmp[8956]*kernel[4]+tmp[8957]*kernel[5]+tmp[9055]*kernel[6]+tmp[9056]*kernel[7]+tmp[9057]*kernel[8];
				ans[8957]<=tmp[8856]*kernel[0]+tmp[8857]*kernel[1]+tmp[8858]*kernel[2]+tmp[8956]*kernel[3]+tmp[8957]*kernel[4]+tmp[8958]*kernel[5]+tmp[9056]*kernel[6]+tmp[9057]*kernel[7]+tmp[9058]*kernel[8];
				ans[8958]<=tmp[8857]*kernel[0]+tmp[8858]*kernel[1]+tmp[8859]*kernel[2]+tmp[8957]*kernel[3]+tmp[8958]*kernel[4]+tmp[8959]*kernel[5]+tmp[9057]*kernel[6]+tmp[9058]*kernel[7]+tmp[9059]*kernel[8];
				ans[8959]<=tmp[8858]*kernel[0]+tmp[8859]*kernel[1]+tmp[8860]*kernel[2]+tmp[8958]*kernel[3]+tmp[8959]*kernel[4]+tmp[8960]*kernel[5]+tmp[9058]*kernel[6]+tmp[9059]*kernel[7]+tmp[9060]*kernel[8];
				ans[8960]<=tmp[8859]*kernel[0]+tmp[8860]*kernel[1]+tmp[8861]*kernel[2]+tmp[8959]*kernel[3]+tmp[8960]*kernel[4]+tmp[8961]*kernel[5]+tmp[9059]*kernel[6]+tmp[9060]*kernel[7]+tmp[9061]*kernel[8];
				ans[8961]<=tmp[8860]*kernel[0]+tmp[8861]*kernel[1]+tmp[8862]*kernel[2]+tmp[8960]*kernel[3]+tmp[8961]*kernel[4]+tmp[8962]*kernel[5]+tmp[9060]*kernel[6]+tmp[9061]*kernel[7]+tmp[9062]*kernel[8];
				ans[8962]<=tmp[8861]*kernel[0]+tmp[8862]*kernel[1]+tmp[8863]*kernel[2]+tmp[8961]*kernel[3]+tmp[8962]*kernel[4]+tmp[8963]*kernel[5]+tmp[9061]*kernel[6]+tmp[9062]*kernel[7]+tmp[9063]*kernel[8];
				ans[8963]<=tmp[8862]*kernel[0]+tmp[8863]*kernel[1]+tmp[8864]*kernel[2]+tmp[8962]*kernel[3]+tmp[8963]*kernel[4]+tmp[8964]*kernel[5]+tmp[9062]*kernel[6]+tmp[9063]*kernel[7]+tmp[9064]*kernel[8];
				ans[8964]<=tmp[8863]*kernel[0]+tmp[8864]*kernel[1]+tmp[8865]*kernel[2]+tmp[8963]*kernel[3]+tmp[8964]*kernel[4]+tmp[8965]*kernel[5]+tmp[9063]*kernel[6]+tmp[9064]*kernel[7]+tmp[9065]*kernel[8];
				ans[8965]<=tmp[8864]*kernel[0]+tmp[8865]*kernel[1]+tmp[8866]*kernel[2]+tmp[8964]*kernel[3]+tmp[8965]*kernel[4]+tmp[8966]*kernel[5]+tmp[9064]*kernel[6]+tmp[9065]*kernel[7]+tmp[9066]*kernel[8];
				ans[8966]<=tmp[8865]*kernel[0]+tmp[8866]*kernel[1]+tmp[8867]*kernel[2]+tmp[8965]*kernel[3]+tmp[8966]*kernel[4]+tmp[8967]*kernel[5]+tmp[9065]*kernel[6]+tmp[9066]*kernel[7]+tmp[9067]*kernel[8];
				ans[8967]<=tmp[8866]*kernel[0]+tmp[8867]*kernel[1]+tmp[8868]*kernel[2]+tmp[8966]*kernel[3]+tmp[8967]*kernel[4]+tmp[8968]*kernel[5]+tmp[9066]*kernel[6]+tmp[9067]*kernel[7]+tmp[9068]*kernel[8];
				ans[8968]<=tmp[8867]*kernel[0]+tmp[8868]*kernel[1]+tmp[8869]*kernel[2]+tmp[8967]*kernel[3]+tmp[8968]*kernel[4]+tmp[8969]*kernel[5]+tmp[9067]*kernel[6]+tmp[9068]*kernel[7]+tmp[9069]*kernel[8];
				ans[8969]<=tmp[8868]*kernel[0]+tmp[8869]*kernel[1]+tmp[8870]*kernel[2]+tmp[8968]*kernel[3]+tmp[8969]*kernel[4]+tmp[8970]*kernel[5]+tmp[9068]*kernel[6]+tmp[9069]*kernel[7]+tmp[9070]*kernel[8];
				ans[8970]<=tmp[8869]*kernel[0]+tmp[8870]*kernel[1]+tmp[8871]*kernel[2]+tmp[8969]*kernel[3]+tmp[8970]*kernel[4]+tmp[8971]*kernel[5]+tmp[9069]*kernel[6]+tmp[9070]*kernel[7]+tmp[9071]*kernel[8];
				ans[8971]<=tmp[8870]*kernel[0]+tmp[8871]*kernel[1]+tmp[8872]*kernel[2]+tmp[8970]*kernel[3]+tmp[8971]*kernel[4]+tmp[8972]*kernel[5]+tmp[9070]*kernel[6]+tmp[9071]*kernel[7]+tmp[9072]*kernel[8];
				ans[8972]<=tmp[8871]*kernel[0]+tmp[8872]*kernel[1]+tmp[8873]*kernel[2]+tmp[8971]*kernel[3]+tmp[8972]*kernel[4]+tmp[8973]*kernel[5]+tmp[9071]*kernel[6]+tmp[9072]*kernel[7]+tmp[9073]*kernel[8];
				ans[8973]<=tmp[8872]*kernel[0]+tmp[8873]*kernel[1]+tmp[8874]*kernel[2]+tmp[8972]*kernel[3]+tmp[8973]*kernel[4]+tmp[8974]*kernel[5]+tmp[9072]*kernel[6]+tmp[9073]*kernel[7]+tmp[9074]*kernel[8];
				ans[8974]<=tmp[8873]*kernel[0]+tmp[8874]*kernel[1]+tmp[8875]*kernel[2]+tmp[8973]*kernel[3]+tmp[8974]*kernel[4]+tmp[8975]*kernel[5]+tmp[9073]*kernel[6]+tmp[9074]*kernel[7]+tmp[9075]*kernel[8];
				ans[8975]<=tmp[8874]*kernel[0]+tmp[8875]*kernel[1]+tmp[8876]*kernel[2]+tmp[8974]*kernel[3]+tmp[8975]*kernel[4]+tmp[8976]*kernel[5]+tmp[9074]*kernel[6]+tmp[9075]*kernel[7]+tmp[9076]*kernel[8];
				ans[8976]<=tmp[8875]*kernel[0]+tmp[8876]*kernel[1]+tmp[8877]*kernel[2]+tmp[8975]*kernel[3]+tmp[8976]*kernel[4]+tmp[8977]*kernel[5]+tmp[9075]*kernel[6]+tmp[9076]*kernel[7]+tmp[9077]*kernel[8];
				ans[8977]<=tmp[8876]*kernel[0]+tmp[8877]*kernel[1]+tmp[8878]*kernel[2]+tmp[8976]*kernel[3]+tmp[8977]*kernel[4]+tmp[8978]*kernel[5]+tmp[9076]*kernel[6]+tmp[9077]*kernel[7]+tmp[9078]*kernel[8];
				ans[8978]<=tmp[8877]*kernel[0]+tmp[8878]*kernel[1]+tmp[8879]*kernel[2]+tmp[8977]*kernel[3]+tmp[8978]*kernel[4]+tmp[8979]*kernel[5]+tmp[9077]*kernel[6]+tmp[9078]*kernel[7]+tmp[9079]*kernel[8];
				ans[8979]<=tmp[8878]*kernel[0]+tmp[8879]*kernel[1]+tmp[8880]*kernel[2]+tmp[8978]*kernel[3]+tmp[8979]*kernel[4]+tmp[8980]*kernel[5]+tmp[9078]*kernel[6]+tmp[9079]*kernel[7]+tmp[9080]*kernel[8];
				ans[8980]<=tmp[8879]*kernel[0]+tmp[8880]*kernel[1]+tmp[8881]*kernel[2]+tmp[8979]*kernel[3]+tmp[8980]*kernel[4]+tmp[8981]*kernel[5]+tmp[9079]*kernel[6]+tmp[9080]*kernel[7]+tmp[9081]*kernel[8];
				ans[8981]<=tmp[8880]*kernel[0]+tmp[8881]*kernel[1]+tmp[8882]*kernel[2]+tmp[8980]*kernel[3]+tmp[8981]*kernel[4]+tmp[8982]*kernel[5]+tmp[9080]*kernel[6]+tmp[9081]*kernel[7]+tmp[9082]*kernel[8];
				ans[8982]<=tmp[8881]*kernel[0]+tmp[8882]*kernel[1]+tmp[8883]*kernel[2]+tmp[8981]*kernel[3]+tmp[8982]*kernel[4]+tmp[8983]*kernel[5]+tmp[9081]*kernel[6]+tmp[9082]*kernel[7]+tmp[9083]*kernel[8];
				ans[8983]<=tmp[8882]*kernel[0]+tmp[8883]*kernel[1]+tmp[8884]*kernel[2]+tmp[8982]*kernel[3]+tmp[8983]*kernel[4]+tmp[8984]*kernel[5]+tmp[9082]*kernel[6]+tmp[9083]*kernel[7]+tmp[9084]*kernel[8];
				ans[8984]<=tmp[8883]*kernel[0]+tmp[8884]*kernel[1]+tmp[8885]*kernel[2]+tmp[8983]*kernel[3]+tmp[8984]*kernel[4]+tmp[8985]*kernel[5]+tmp[9083]*kernel[6]+tmp[9084]*kernel[7]+tmp[9085]*kernel[8];
				ans[8985]<=tmp[8884]*kernel[0]+tmp[8885]*kernel[1]+tmp[8886]*kernel[2]+tmp[8984]*kernel[3]+tmp[8985]*kernel[4]+tmp[8986]*kernel[5]+tmp[9084]*kernel[6]+tmp[9085]*kernel[7]+tmp[9086]*kernel[8];
				ans[8986]<=tmp[8885]*kernel[0]+tmp[8886]*kernel[1]+tmp[8887]*kernel[2]+tmp[8985]*kernel[3]+tmp[8986]*kernel[4]+tmp[8987]*kernel[5]+tmp[9085]*kernel[6]+tmp[9086]*kernel[7]+tmp[9087]*kernel[8];
				ans[8987]<=tmp[8886]*kernel[0]+tmp[8887]*kernel[1]+tmp[8888]*kernel[2]+tmp[8986]*kernel[3]+tmp[8987]*kernel[4]+tmp[8988]*kernel[5]+tmp[9086]*kernel[6]+tmp[9087]*kernel[7]+tmp[9088]*kernel[8];
				ans[8988]<=tmp[8887]*kernel[0]+tmp[8888]*kernel[1]+tmp[8889]*kernel[2]+tmp[8987]*kernel[3]+tmp[8988]*kernel[4]+tmp[8989]*kernel[5]+tmp[9087]*kernel[6]+tmp[9088]*kernel[7]+tmp[9089]*kernel[8];
				ans[8989]<=tmp[8888]*kernel[0]+tmp[8889]*kernel[1]+tmp[8890]*kernel[2]+tmp[8988]*kernel[3]+tmp[8989]*kernel[4]+tmp[8990]*kernel[5]+tmp[9088]*kernel[6]+tmp[9089]*kernel[7]+tmp[9090]*kernel[8];
				ans[8990]<=tmp[8889]*kernel[0]+tmp[8890]*kernel[1]+tmp[8891]*kernel[2]+tmp[8989]*kernel[3]+tmp[8990]*kernel[4]+tmp[8991]*kernel[5]+tmp[9089]*kernel[6]+tmp[9090]*kernel[7]+tmp[9091]*kernel[8];
				ans[8991]<=tmp[8890]*kernel[0]+tmp[8891]*kernel[1]+tmp[8892]*kernel[2]+tmp[8990]*kernel[3]+tmp[8991]*kernel[4]+tmp[8992]*kernel[5]+tmp[9090]*kernel[6]+tmp[9091]*kernel[7]+tmp[9092]*kernel[8];
				ans[8992]<=tmp[8891]*kernel[0]+tmp[8892]*kernel[1]+tmp[8893]*kernel[2]+tmp[8991]*kernel[3]+tmp[8992]*kernel[4]+tmp[8993]*kernel[5]+tmp[9091]*kernel[6]+tmp[9092]*kernel[7]+tmp[9093]*kernel[8];
				ans[8993]<=tmp[8892]*kernel[0]+tmp[8893]*kernel[1]+tmp[8894]*kernel[2]+tmp[8992]*kernel[3]+tmp[8993]*kernel[4]+tmp[8994]*kernel[5]+tmp[9092]*kernel[6]+tmp[9093]*kernel[7]+tmp[9094]*kernel[8];
				ans[8994]<=tmp[8893]*kernel[0]+tmp[8894]*kernel[1]+tmp[8895]*kernel[2]+tmp[8993]*kernel[3]+tmp[8994]*kernel[4]+tmp[8995]*kernel[5]+tmp[9093]*kernel[6]+tmp[9094]*kernel[7]+tmp[9095]*kernel[8];
				ans[8995]<=tmp[8894]*kernel[0]+tmp[8895]*kernel[1]+tmp[8896]*kernel[2]+tmp[8994]*kernel[3]+tmp[8995]*kernel[4]+tmp[8996]*kernel[5]+tmp[9094]*kernel[6]+tmp[9095]*kernel[7]+tmp[9096]*kernel[8];
				ans[8996]<=tmp[8895]*kernel[0]+tmp[8896]*kernel[1]+tmp[8897]*kernel[2]+tmp[8995]*kernel[3]+tmp[8996]*kernel[4]+tmp[8997]*kernel[5]+tmp[9095]*kernel[6]+tmp[9096]*kernel[7]+tmp[9097]*kernel[8];
				ans[8997]<=tmp[8896]*kernel[0]+tmp[8897]*kernel[1]+tmp[8898]*kernel[2]+tmp[8996]*kernel[3]+tmp[8997]*kernel[4]+tmp[8998]*kernel[5]+tmp[9096]*kernel[6]+tmp[9097]*kernel[7]+tmp[9098]*kernel[8];
				ans[8998]<=tmp[8897]*kernel[0]+tmp[8898]*kernel[1]+tmp[8899]*kernel[2]+tmp[8997]*kernel[3]+tmp[8998]*kernel[4]+tmp[8999]*kernel[5]+tmp[9097]*kernel[6]+tmp[9098]*kernel[7]+tmp[9099]*kernel[8];
				ans[8999]<=tmp[8898]*kernel[0]+tmp[8899]*kernel[1]+tmp[8998]*kernel[3]+tmp[8999]*kernel[4]+tmp[9098]*kernel[6]+tmp[9099]*kernel[7];
				ans[9000]<=tmp[8900]*kernel[1]+tmp[8901]*kernel[2]+tmp[9000]*kernel[4]+tmp[9001]*kernel[5]+tmp[9100]*kernel[7]+tmp[9101]*kernel[8];
				ans[9001]<=tmp[8900]*kernel[0]+tmp[8901]*kernel[1]+tmp[8902]*kernel[2]+tmp[9000]*kernel[3]+tmp[9001]*kernel[4]+tmp[9002]*kernel[5]+tmp[9100]*kernel[6]+tmp[9101]*kernel[7]+tmp[9102]*kernel[8];
				ans[9002]<=tmp[8901]*kernel[0]+tmp[8902]*kernel[1]+tmp[8903]*kernel[2]+tmp[9001]*kernel[3]+tmp[9002]*kernel[4]+tmp[9003]*kernel[5]+tmp[9101]*kernel[6]+tmp[9102]*kernel[7]+tmp[9103]*kernel[8];
				ans[9003]<=tmp[8902]*kernel[0]+tmp[8903]*kernel[1]+tmp[8904]*kernel[2]+tmp[9002]*kernel[3]+tmp[9003]*kernel[4]+tmp[9004]*kernel[5]+tmp[9102]*kernel[6]+tmp[9103]*kernel[7]+tmp[9104]*kernel[8];
				ans[9004]<=tmp[8903]*kernel[0]+tmp[8904]*kernel[1]+tmp[8905]*kernel[2]+tmp[9003]*kernel[3]+tmp[9004]*kernel[4]+tmp[9005]*kernel[5]+tmp[9103]*kernel[6]+tmp[9104]*kernel[7]+tmp[9105]*kernel[8];
				ans[9005]<=tmp[8904]*kernel[0]+tmp[8905]*kernel[1]+tmp[8906]*kernel[2]+tmp[9004]*kernel[3]+tmp[9005]*kernel[4]+tmp[9006]*kernel[5]+tmp[9104]*kernel[6]+tmp[9105]*kernel[7]+tmp[9106]*kernel[8];
				ans[9006]<=tmp[8905]*kernel[0]+tmp[8906]*kernel[1]+tmp[8907]*kernel[2]+tmp[9005]*kernel[3]+tmp[9006]*kernel[4]+tmp[9007]*kernel[5]+tmp[9105]*kernel[6]+tmp[9106]*kernel[7]+tmp[9107]*kernel[8];
				ans[9007]<=tmp[8906]*kernel[0]+tmp[8907]*kernel[1]+tmp[8908]*kernel[2]+tmp[9006]*kernel[3]+tmp[9007]*kernel[4]+tmp[9008]*kernel[5]+tmp[9106]*kernel[6]+tmp[9107]*kernel[7]+tmp[9108]*kernel[8];
				ans[9008]<=tmp[8907]*kernel[0]+tmp[8908]*kernel[1]+tmp[8909]*kernel[2]+tmp[9007]*kernel[3]+tmp[9008]*kernel[4]+tmp[9009]*kernel[5]+tmp[9107]*kernel[6]+tmp[9108]*kernel[7]+tmp[9109]*kernel[8];
				ans[9009]<=tmp[8908]*kernel[0]+tmp[8909]*kernel[1]+tmp[8910]*kernel[2]+tmp[9008]*kernel[3]+tmp[9009]*kernel[4]+tmp[9010]*kernel[5]+tmp[9108]*kernel[6]+tmp[9109]*kernel[7]+tmp[9110]*kernel[8];
				ans[9010]<=tmp[8909]*kernel[0]+tmp[8910]*kernel[1]+tmp[8911]*kernel[2]+tmp[9009]*kernel[3]+tmp[9010]*kernel[4]+tmp[9011]*kernel[5]+tmp[9109]*kernel[6]+tmp[9110]*kernel[7]+tmp[9111]*kernel[8];
				ans[9011]<=tmp[8910]*kernel[0]+tmp[8911]*kernel[1]+tmp[8912]*kernel[2]+tmp[9010]*kernel[3]+tmp[9011]*kernel[4]+tmp[9012]*kernel[5]+tmp[9110]*kernel[6]+tmp[9111]*kernel[7]+tmp[9112]*kernel[8];
				ans[9012]<=tmp[8911]*kernel[0]+tmp[8912]*kernel[1]+tmp[8913]*kernel[2]+tmp[9011]*kernel[3]+tmp[9012]*kernel[4]+tmp[9013]*kernel[5]+tmp[9111]*kernel[6]+tmp[9112]*kernel[7]+tmp[9113]*kernel[8];
				ans[9013]<=tmp[8912]*kernel[0]+tmp[8913]*kernel[1]+tmp[8914]*kernel[2]+tmp[9012]*kernel[3]+tmp[9013]*kernel[4]+tmp[9014]*kernel[5]+tmp[9112]*kernel[6]+tmp[9113]*kernel[7]+tmp[9114]*kernel[8];
				ans[9014]<=tmp[8913]*kernel[0]+tmp[8914]*kernel[1]+tmp[8915]*kernel[2]+tmp[9013]*kernel[3]+tmp[9014]*kernel[4]+tmp[9015]*kernel[5]+tmp[9113]*kernel[6]+tmp[9114]*kernel[7]+tmp[9115]*kernel[8];
				ans[9015]<=tmp[8914]*kernel[0]+tmp[8915]*kernel[1]+tmp[8916]*kernel[2]+tmp[9014]*kernel[3]+tmp[9015]*kernel[4]+tmp[9016]*kernel[5]+tmp[9114]*kernel[6]+tmp[9115]*kernel[7]+tmp[9116]*kernel[8];
				ans[9016]<=tmp[8915]*kernel[0]+tmp[8916]*kernel[1]+tmp[8917]*kernel[2]+tmp[9015]*kernel[3]+tmp[9016]*kernel[4]+tmp[9017]*kernel[5]+tmp[9115]*kernel[6]+tmp[9116]*kernel[7]+tmp[9117]*kernel[8];
				ans[9017]<=tmp[8916]*kernel[0]+tmp[8917]*kernel[1]+tmp[8918]*kernel[2]+tmp[9016]*kernel[3]+tmp[9017]*kernel[4]+tmp[9018]*kernel[5]+tmp[9116]*kernel[6]+tmp[9117]*kernel[7]+tmp[9118]*kernel[8];
				ans[9018]<=tmp[8917]*kernel[0]+tmp[8918]*kernel[1]+tmp[8919]*kernel[2]+tmp[9017]*kernel[3]+tmp[9018]*kernel[4]+tmp[9019]*kernel[5]+tmp[9117]*kernel[6]+tmp[9118]*kernel[7]+tmp[9119]*kernel[8];
				ans[9019]<=tmp[8918]*kernel[0]+tmp[8919]*kernel[1]+tmp[8920]*kernel[2]+tmp[9018]*kernel[3]+tmp[9019]*kernel[4]+tmp[9020]*kernel[5]+tmp[9118]*kernel[6]+tmp[9119]*kernel[7]+tmp[9120]*kernel[8];
				ans[9020]<=tmp[8919]*kernel[0]+tmp[8920]*kernel[1]+tmp[8921]*kernel[2]+tmp[9019]*kernel[3]+tmp[9020]*kernel[4]+tmp[9021]*kernel[5]+tmp[9119]*kernel[6]+tmp[9120]*kernel[7]+tmp[9121]*kernel[8];
				ans[9021]<=tmp[8920]*kernel[0]+tmp[8921]*kernel[1]+tmp[8922]*kernel[2]+tmp[9020]*kernel[3]+tmp[9021]*kernel[4]+tmp[9022]*kernel[5]+tmp[9120]*kernel[6]+tmp[9121]*kernel[7]+tmp[9122]*kernel[8];
				ans[9022]<=tmp[8921]*kernel[0]+tmp[8922]*kernel[1]+tmp[8923]*kernel[2]+tmp[9021]*kernel[3]+tmp[9022]*kernel[4]+tmp[9023]*kernel[5]+tmp[9121]*kernel[6]+tmp[9122]*kernel[7]+tmp[9123]*kernel[8];
				ans[9023]<=tmp[8922]*kernel[0]+tmp[8923]*kernel[1]+tmp[8924]*kernel[2]+tmp[9022]*kernel[3]+tmp[9023]*kernel[4]+tmp[9024]*kernel[5]+tmp[9122]*kernel[6]+tmp[9123]*kernel[7]+tmp[9124]*kernel[8];
				ans[9024]<=tmp[8923]*kernel[0]+tmp[8924]*kernel[1]+tmp[8925]*kernel[2]+tmp[9023]*kernel[3]+tmp[9024]*kernel[4]+tmp[9025]*kernel[5]+tmp[9123]*kernel[6]+tmp[9124]*kernel[7]+tmp[9125]*kernel[8];
				ans[9025]<=tmp[8924]*kernel[0]+tmp[8925]*kernel[1]+tmp[8926]*kernel[2]+tmp[9024]*kernel[3]+tmp[9025]*kernel[4]+tmp[9026]*kernel[5]+tmp[9124]*kernel[6]+tmp[9125]*kernel[7]+tmp[9126]*kernel[8];
				ans[9026]<=tmp[8925]*kernel[0]+tmp[8926]*kernel[1]+tmp[8927]*kernel[2]+tmp[9025]*kernel[3]+tmp[9026]*kernel[4]+tmp[9027]*kernel[5]+tmp[9125]*kernel[6]+tmp[9126]*kernel[7]+tmp[9127]*kernel[8];
				ans[9027]<=tmp[8926]*kernel[0]+tmp[8927]*kernel[1]+tmp[8928]*kernel[2]+tmp[9026]*kernel[3]+tmp[9027]*kernel[4]+tmp[9028]*kernel[5]+tmp[9126]*kernel[6]+tmp[9127]*kernel[7]+tmp[9128]*kernel[8];
				ans[9028]<=tmp[8927]*kernel[0]+tmp[8928]*kernel[1]+tmp[8929]*kernel[2]+tmp[9027]*kernel[3]+tmp[9028]*kernel[4]+tmp[9029]*kernel[5]+tmp[9127]*kernel[6]+tmp[9128]*kernel[7]+tmp[9129]*kernel[8];
				ans[9029]<=tmp[8928]*kernel[0]+tmp[8929]*kernel[1]+tmp[8930]*kernel[2]+tmp[9028]*kernel[3]+tmp[9029]*kernel[4]+tmp[9030]*kernel[5]+tmp[9128]*kernel[6]+tmp[9129]*kernel[7]+tmp[9130]*kernel[8];
				ans[9030]<=tmp[8929]*kernel[0]+tmp[8930]*kernel[1]+tmp[8931]*kernel[2]+tmp[9029]*kernel[3]+tmp[9030]*kernel[4]+tmp[9031]*kernel[5]+tmp[9129]*kernel[6]+tmp[9130]*kernel[7]+tmp[9131]*kernel[8];
				ans[9031]<=tmp[8930]*kernel[0]+tmp[8931]*kernel[1]+tmp[8932]*kernel[2]+tmp[9030]*kernel[3]+tmp[9031]*kernel[4]+tmp[9032]*kernel[5]+tmp[9130]*kernel[6]+tmp[9131]*kernel[7]+tmp[9132]*kernel[8];
				ans[9032]<=tmp[8931]*kernel[0]+tmp[8932]*kernel[1]+tmp[8933]*kernel[2]+tmp[9031]*kernel[3]+tmp[9032]*kernel[4]+tmp[9033]*kernel[5]+tmp[9131]*kernel[6]+tmp[9132]*kernel[7]+tmp[9133]*kernel[8];
				ans[9033]<=tmp[8932]*kernel[0]+tmp[8933]*kernel[1]+tmp[8934]*kernel[2]+tmp[9032]*kernel[3]+tmp[9033]*kernel[4]+tmp[9034]*kernel[5]+tmp[9132]*kernel[6]+tmp[9133]*kernel[7]+tmp[9134]*kernel[8];
				ans[9034]<=tmp[8933]*kernel[0]+tmp[8934]*kernel[1]+tmp[8935]*kernel[2]+tmp[9033]*kernel[3]+tmp[9034]*kernel[4]+tmp[9035]*kernel[5]+tmp[9133]*kernel[6]+tmp[9134]*kernel[7]+tmp[9135]*kernel[8];
				ans[9035]<=tmp[8934]*kernel[0]+tmp[8935]*kernel[1]+tmp[8936]*kernel[2]+tmp[9034]*kernel[3]+tmp[9035]*kernel[4]+tmp[9036]*kernel[5]+tmp[9134]*kernel[6]+tmp[9135]*kernel[7]+tmp[9136]*kernel[8];
				ans[9036]<=tmp[8935]*kernel[0]+tmp[8936]*kernel[1]+tmp[8937]*kernel[2]+tmp[9035]*kernel[3]+tmp[9036]*kernel[4]+tmp[9037]*kernel[5]+tmp[9135]*kernel[6]+tmp[9136]*kernel[7]+tmp[9137]*kernel[8];
				ans[9037]<=tmp[8936]*kernel[0]+tmp[8937]*kernel[1]+tmp[8938]*kernel[2]+tmp[9036]*kernel[3]+tmp[9037]*kernel[4]+tmp[9038]*kernel[5]+tmp[9136]*kernel[6]+tmp[9137]*kernel[7]+tmp[9138]*kernel[8];
				ans[9038]<=tmp[8937]*kernel[0]+tmp[8938]*kernel[1]+tmp[8939]*kernel[2]+tmp[9037]*kernel[3]+tmp[9038]*kernel[4]+tmp[9039]*kernel[5]+tmp[9137]*kernel[6]+tmp[9138]*kernel[7]+tmp[9139]*kernel[8];
				ans[9039]<=tmp[8938]*kernel[0]+tmp[8939]*kernel[1]+tmp[8940]*kernel[2]+tmp[9038]*kernel[3]+tmp[9039]*kernel[4]+tmp[9040]*kernel[5]+tmp[9138]*kernel[6]+tmp[9139]*kernel[7]+tmp[9140]*kernel[8];
				ans[9040]<=tmp[8939]*kernel[0]+tmp[8940]*kernel[1]+tmp[8941]*kernel[2]+tmp[9039]*kernel[3]+tmp[9040]*kernel[4]+tmp[9041]*kernel[5]+tmp[9139]*kernel[6]+tmp[9140]*kernel[7]+tmp[9141]*kernel[8];
				ans[9041]<=tmp[8940]*kernel[0]+tmp[8941]*kernel[1]+tmp[8942]*kernel[2]+tmp[9040]*kernel[3]+tmp[9041]*kernel[4]+tmp[9042]*kernel[5]+tmp[9140]*kernel[6]+tmp[9141]*kernel[7]+tmp[9142]*kernel[8];
				ans[9042]<=tmp[8941]*kernel[0]+tmp[8942]*kernel[1]+tmp[8943]*kernel[2]+tmp[9041]*kernel[3]+tmp[9042]*kernel[4]+tmp[9043]*kernel[5]+tmp[9141]*kernel[6]+tmp[9142]*kernel[7]+tmp[9143]*kernel[8];
				ans[9043]<=tmp[8942]*kernel[0]+tmp[8943]*kernel[1]+tmp[8944]*kernel[2]+tmp[9042]*kernel[3]+tmp[9043]*kernel[4]+tmp[9044]*kernel[5]+tmp[9142]*kernel[6]+tmp[9143]*kernel[7]+tmp[9144]*kernel[8];
				ans[9044]<=tmp[8943]*kernel[0]+tmp[8944]*kernel[1]+tmp[8945]*kernel[2]+tmp[9043]*kernel[3]+tmp[9044]*kernel[4]+tmp[9045]*kernel[5]+tmp[9143]*kernel[6]+tmp[9144]*kernel[7]+tmp[9145]*kernel[8];
				ans[9045]<=tmp[8944]*kernel[0]+tmp[8945]*kernel[1]+tmp[8946]*kernel[2]+tmp[9044]*kernel[3]+tmp[9045]*kernel[4]+tmp[9046]*kernel[5]+tmp[9144]*kernel[6]+tmp[9145]*kernel[7]+tmp[9146]*kernel[8];
				ans[9046]<=tmp[8945]*kernel[0]+tmp[8946]*kernel[1]+tmp[8947]*kernel[2]+tmp[9045]*kernel[3]+tmp[9046]*kernel[4]+tmp[9047]*kernel[5]+tmp[9145]*kernel[6]+tmp[9146]*kernel[7]+tmp[9147]*kernel[8];
				ans[9047]<=tmp[8946]*kernel[0]+tmp[8947]*kernel[1]+tmp[8948]*kernel[2]+tmp[9046]*kernel[3]+tmp[9047]*kernel[4]+tmp[9048]*kernel[5]+tmp[9146]*kernel[6]+tmp[9147]*kernel[7]+tmp[9148]*kernel[8];
				ans[9048]<=tmp[8947]*kernel[0]+tmp[8948]*kernel[1]+tmp[8949]*kernel[2]+tmp[9047]*kernel[3]+tmp[9048]*kernel[4]+tmp[9049]*kernel[5]+tmp[9147]*kernel[6]+tmp[9148]*kernel[7]+tmp[9149]*kernel[8];
				ans[9049]<=tmp[8948]*kernel[0]+tmp[8949]*kernel[1]+tmp[8950]*kernel[2]+tmp[9048]*kernel[3]+tmp[9049]*kernel[4]+tmp[9050]*kernel[5]+tmp[9148]*kernel[6]+tmp[9149]*kernel[7]+tmp[9150]*kernel[8];
				ans[9050]<=tmp[8949]*kernel[0]+tmp[8950]*kernel[1]+tmp[8951]*kernel[2]+tmp[9049]*kernel[3]+tmp[9050]*kernel[4]+tmp[9051]*kernel[5]+tmp[9149]*kernel[6]+tmp[9150]*kernel[7]+tmp[9151]*kernel[8];
				ans[9051]<=tmp[8950]*kernel[0]+tmp[8951]*kernel[1]+tmp[8952]*kernel[2]+tmp[9050]*kernel[3]+tmp[9051]*kernel[4]+tmp[9052]*kernel[5]+tmp[9150]*kernel[6]+tmp[9151]*kernel[7]+tmp[9152]*kernel[8];
				ans[9052]<=tmp[8951]*kernel[0]+tmp[8952]*kernel[1]+tmp[8953]*kernel[2]+tmp[9051]*kernel[3]+tmp[9052]*kernel[4]+tmp[9053]*kernel[5]+tmp[9151]*kernel[6]+tmp[9152]*kernel[7]+tmp[9153]*kernel[8];
				ans[9053]<=tmp[8952]*kernel[0]+tmp[8953]*kernel[1]+tmp[8954]*kernel[2]+tmp[9052]*kernel[3]+tmp[9053]*kernel[4]+tmp[9054]*kernel[5]+tmp[9152]*kernel[6]+tmp[9153]*kernel[7]+tmp[9154]*kernel[8];
				ans[9054]<=tmp[8953]*kernel[0]+tmp[8954]*kernel[1]+tmp[8955]*kernel[2]+tmp[9053]*kernel[3]+tmp[9054]*kernel[4]+tmp[9055]*kernel[5]+tmp[9153]*kernel[6]+tmp[9154]*kernel[7]+tmp[9155]*kernel[8];
				ans[9055]<=tmp[8954]*kernel[0]+tmp[8955]*kernel[1]+tmp[8956]*kernel[2]+tmp[9054]*kernel[3]+tmp[9055]*kernel[4]+tmp[9056]*kernel[5]+tmp[9154]*kernel[6]+tmp[9155]*kernel[7]+tmp[9156]*kernel[8];
				ans[9056]<=tmp[8955]*kernel[0]+tmp[8956]*kernel[1]+tmp[8957]*kernel[2]+tmp[9055]*kernel[3]+tmp[9056]*kernel[4]+tmp[9057]*kernel[5]+tmp[9155]*kernel[6]+tmp[9156]*kernel[7]+tmp[9157]*kernel[8];
				ans[9057]<=tmp[8956]*kernel[0]+tmp[8957]*kernel[1]+tmp[8958]*kernel[2]+tmp[9056]*kernel[3]+tmp[9057]*kernel[4]+tmp[9058]*kernel[5]+tmp[9156]*kernel[6]+tmp[9157]*kernel[7]+tmp[9158]*kernel[8];
				ans[9058]<=tmp[8957]*kernel[0]+tmp[8958]*kernel[1]+tmp[8959]*kernel[2]+tmp[9057]*kernel[3]+tmp[9058]*kernel[4]+tmp[9059]*kernel[5]+tmp[9157]*kernel[6]+tmp[9158]*kernel[7]+tmp[9159]*kernel[8];
				ans[9059]<=tmp[8958]*kernel[0]+tmp[8959]*kernel[1]+tmp[8960]*kernel[2]+tmp[9058]*kernel[3]+tmp[9059]*kernel[4]+tmp[9060]*kernel[5]+tmp[9158]*kernel[6]+tmp[9159]*kernel[7]+tmp[9160]*kernel[8];
				ans[9060]<=tmp[8959]*kernel[0]+tmp[8960]*kernel[1]+tmp[8961]*kernel[2]+tmp[9059]*kernel[3]+tmp[9060]*kernel[4]+tmp[9061]*kernel[5]+tmp[9159]*kernel[6]+tmp[9160]*kernel[7]+tmp[9161]*kernel[8];
				ans[9061]<=tmp[8960]*kernel[0]+tmp[8961]*kernel[1]+tmp[8962]*kernel[2]+tmp[9060]*kernel[3]+tmp[9061]*kernel[4]+tmp[9062]*kernel[5]+tmp[9160]*kernel[6]+tmp[9161]*kernel[7]+tmp[9162]*kernel[8];
				ans[9062]<=tmp[8961]*kernel[0]+tmp[8962]*kernel[1]+tmp[8963]*kernel[2]+tmp[9061]*kernel[3]+tmp[9062]*kernel[4]+tmp[9063]*kernel[5]+tmp[9161]*kernel[6]+tmp[9162]*kernel[7]+tmp[9163]*kernel[8];
				ans[9063]<=tmp[8962]*kernel[0]+tmp[8963]*kernel[1]+tmp[8964]*kernel[2]+tmp[9062]*kernel[3]+tmp[9063]*kernel[4]+tmp[9064]*kernel[5]+tmp[9162]*kernel[6]+tmp[9163]*kernel[7]+tmp[9164]*kernel[8];
				ans[9064]<=tmp[8963]*kernel[0]+tmp[8964]*kernel[1]+tmp[8965]*kernel[2]+tmp[9063]*kernel[3]+tmp[9064]*kernel[4]+tmp[9065]*kernel[5]+tmp[9163]*kernel[6]+tmp[9164]*kernel[7]+tmp[9165]*kernel[8];
				ans[9065]<=tmp[8964]*kernel[0]+tmp[8965]*kernel[1]+tmp[8966]*kernel[2]+tmp[9064]*kernel[3]+tmp[9065]*kernel[4]+tmp[9066]*kernel[5]+tmp[9164]*kernel[6]+tmp[9165]*kernel[7]+tmp[9166]*kernel[8];
				ans[9066]<=tmp[8965]*kernel[0]+tmp[8966]*kernel[1]+tmp[8967]*kernel[2]+tmp[9065]*kernel[3]+tmp[9066]*kernel[4]+tmp[9067]*kernel[5]+tmp[9165]*kernel[6]+tmp[9166]*kernel[7]+tmp[9167]*kernel[8];
				ans[9067]<=tmp[8966]*kernel[0]+tmp[8967]*kernel[1]+tmp[8968]*kernel[2]+tmp[9066]*kernel[3]+tmp[9067]*kernel[4]+tmp[9068]*kernel[5]+tmp[9166]*kernel[6]+tmp[9167]*kernel[7]+tmp[9168]*kernel[8];
				ans[9068]<=tmp[8967]*kernel[0]+tmp[8968]*kernel[1]+tmp[8969]*kernel[2]+tmp[9067]*kernel[3]+tmp[9068]*kernel[4]+tmp[9069]*kernel[5]+tmp[9167]*kernel[6]+tmp[9168]*kernel[7]+tmp[9169]*kernel[8];
				ans[9069]<=tmp[8968]*kernel[0]+tmp[8969]*kernel[1]+tmp[8970]*kernel[2]+tmp[9068]*kernel[3]+tmp[9069]*kernel[4]+tmp[9070]*kernel[5]+tmp[9168]*kernel[6]+tmp[9169]*kernel[7]+tmp[9170]*kernel[8];
				ans[9070]<=tmp[8969]*kernel[0]+tmp[8970]*kernel[1]+tmp[8971]*kernel[2]+tmp[9069]*kernel[3]+tmp[9070]*kernel[4]+tmp[9071]*kernel[5]+tmp[9169]*kernel[6]+tmp[9170]*kernel[7]+tmp[9171]*kernel[8];
				ans[9071]<=tmp[8970]*kernel[0]+tmp[8971]*kernel[1]+tmp[8972]*kernel[2]+tmp[9070]*kernel[3]+tmp[9071]*kernel[4]+tmp[9072]*kernel[5]+tmp[9170]*kernel[6]+tmp[9171]*kernel[7]+tmp[9172]*kernel[8];
				ans[9072]<=tmp[8971]*kernel[0]+tmp[8972]*kernel[1]+tmp[8973]*kernel[2]+tmp[9071]*kernel[3]+tmp[9072]*kernel[4]+tmp[9073]*kernel[5]+tmp[9171]*kernel[6]+tmp[9172]*kernel[7]+tmp[9173]*kernel[8];
				ans[9073]<=tmp[8972]*kernel[0]+tmp[8973]*kernel[1]+tmp[8974]*kernel[2]+tmp[9072]*kernel[3]+tmp[9073]*kernel[4]+tmp[9074]*kernel[5]+tmp[9172]*kernel[6]+tmp[9173]*kernel[7]+tmp[9174]*kernel[8];
				ans[9074]<=tmp[8973]*kernel[0]+tmp[8974]*kernel[1]+tmp[8975]*kernel[2]+tmp[9073]*kernel[3]+tmp[9074]*kernel[4]+tmp[9075]*kernel[5]+tmp[9173]*kernel[6]+tmp[9174]*kernel[7]+tmp[9175]*kernel[8];
				ans[9075]<=tmp[8974]*kernel[0]+tmp[8975]*kernel[1]+tmp[8976]*kernel[2]+tmp[9074]*kernel[3]+tmp[9075]*kernel[4]+tmp[9076]*kernel[5]+tmp[9174]*kernel[6]+tmp[9175]*kernel[7]+tmp[9176]*kernel[8];
				ans[9076]<=tmp[8975]*kernel[0]+tmp[8976]*kernel[1]+tmp[8977]*kernel[2]+tmp[9075]*kernel[3]+tmp[9076]*kernel[4]+tmp[9077]*kernel[5]+tmp[9175]*kernel[6]+tmp[9176]*kernel[7]+tmp[9177]*kernel[8];
				ans[9077]<=tmp[8976]*kernel[0]+tmp[8977]*kernel[1]+tmp[8978]*kernel[2]+tmp[9076]*kernel[3]+tmp[9077]*kernel[4]+tmp[9078]*kernel[5]+tmp[9176]*kernel[6]+tmp[9177]*kernel[7]+tmp[9178]*kernel[8];
				ans[9078]<=tmp[8977]*kernel[0]+tmp[8978]*kernel[1]+tmp[8979]*kernel[2]+tmp[9077]*kernel[3]+tmp[9078]*kernel[4]+tmp[9079]*kernel[5]+tmp[9177]*kernel[6]+tmp[9178]*kernel[7]+tmp[9179]*kernel[8];
				ans[9079]<=tmp[8978]*kernel[0]+tmp[8979]*kernel[1]+tmp[8980]*kernel[2]+tmp[9078]*kernel[3]+tmp[9079]*kernel[4]+tmp[9080]*kernel[5]+tmp[9178]*kernel[6]+tmp[9179]*kernel[7]+tmp[9180]*kernel[8];
				ans[9080]<=tmp[8979]*kernel[0]+tmp[8980]*kernel[1]+tmp[8981]*kernel[2]+tmp[9079]*kernel[3]+tmp[9080]*kernel[4]+tmp[9081]*kernel[5]+tmp[9179]*kernel[6]+tmp[9180]*kernel[7]+tmp[9181]*kernel[8];
				ans[9081]<=tmp[8980]*kernel[0]+tmp[8981]*kernel[1]+tmp[8982]*kernel[2]+tmp[9080]*kernel[3]+tmp[9081]*kernel[4]+tmp[9082]*kernel[5]+tmp[9180]*kernel[6]+tmp[9181]*kernel[7]+tmp[9182]*kernel[8];
				ans[9082]<=tmp[8981]*kernel[0]+tmp[8982]*kernel[1]+tmp[8983]*kernel[2]+tmp[9081]*kernel[3]+tmp[9082]*kernel[4]+tmp[9083]*kernel[5]+tmp[9181]*kernel[6]+tmp[9182]*kernel[7]+tmp[9183]*kernel[8];
				ans[9083]<=tmp[8982]*kernel[0]+tmp[8983]*kernel[1]+tmp[8984]*kernel[2]+tmp[9082]*kernel[3]+tmp[9083]*kernel[4]+tmp[9084]*kernel[5]+tmp[9182]*kernel[6]+tmp[9183]*kernel[7]+tmp[9184]*kernel[8];
				ans[9084]<=tmp[8983]*kernel[0]+tmp[8984]*kernel[1]+tmp[8985]*kernel[2]+tmp[9083]*kernel[3]+tmp[9084]*kernel[4]+tmp[9085]*kernel[5]+tmp[9183]*kernel[6]+tmp[9184]*kernel[7]+tmp[9185]*kernel[8];
				ans[9085]<=tmp[8984]*kernel[0]+tmp[8985]*kernel[1]+tmp[8986]*kernel[2]+tmp[9084]*kernel[3]+tmp[9085]*kernel[4]+tmp[9086]*kernel[5]+tmp[9184]*kernel[6]+tmp[9185]*kernel[7]+tmp[9186]*kernel[8];
				ans[9086]<=tmp[8985]*kernel[0]+tmp[8986]*kernel[1]+tmp[8987]*kernel[2]+tmp[9085]*kernel[3]+tmp[9086]*kernel[4]+tmp[9087]*kernel[5]+tmp[9185]*kernel[6]+tmp[9186]*kernel[7]+tmp[9187]*kernel[8];
				ans[9087]<=tmp[8986]*kernel[0]+tmp[8987]*kernel[1]+tmp[8988]*kernel[2]+tmp[9086]*kernel[3]+tmp[9087]*kernel[4]+tmp[9088]*kernel[5]+tmp[9186]*kernel[6]+tmp[9187]*kernel[7]+tmp[9188]*kernel[8];
				ans[9088]<=tmp[8987]*kernel[0]+tmp[8988]*kernel[1]+tmp[8989]*kernel[2]+tmp[9087]*kernel[3]+tmp[9088]*kernel[4]+tmp[9089]*kernel[5]+tmp[9187]*kernel[6]+tmp[9188]*kernel[7]+tmp[9189]*kernel[8];
				ans[9089]<=tmp[8988]*kernel[0]+tmp[8989]*kernel[1]+tmp[8990]*kernel[2]+tmp[9088]*kernel[3]+tmp[9089]*kernel[4]+tmp[9090]*kernel[5]+tmp[9188]*kernel[6]+tmp[9189]*kernel[7]+tmp[9190]*kernel[8];
				ans[9090]<=tmp[8989]*kernel[0]+tmp[8990]*kernel[1]+tmp[8991]*kernel[2]+tmp[9089]*kernel[3]+tmp[9090]*kernel[4]+tmp[9091]*kernel[5]+tmp[9189]*kernel[6]+tmp[9190]*kernel[7]+tmp[9191]*kernel[8];
				ans[9091]<=tmp[8990]*kernel[0]+tmp[8991]*kernel[1]+tmp[8992]*kernel[2]+tmp[9090]*kernel[3]+tmp[9091]*kernel[4]+tmp[9092]*kernel[5]+tmp[9190]*kernel[6]+tmp[9191]*kernel[7]+tmp[9192]*kernel[8];
				ans[9092]<=tmp[8991]*kernel[0]+tmp[8992]*kernel[1]+tmp[8993]*kernel[2]+tmp[9091]*kernel[3]+tmp[9092]*kernel[4]+tmp[9093]*kernel[5]+tmp[9191]*kernel[6]+tmp[9192]*kernel[7]+tmp[9193]*kernel[8];
				ans[9093]<=tmp[8992]*kernel[0]+tmp[8993]*kernel[1]+tmp[8994]*kernel[2]+tmp[9092]*kernel[3]+tmp[9093]*kernel[4]+tmp[9094]*kernel[5]+tmp[9192]*kernel[6]+tmp[9193]*kernel[7]+tmp[9194]*kernel[8];
				ans[9094]<=tmp[8993]*kernel[0]+tmp[8994]*kernel[1]+tmp[8995]*kernel[2]+tmp[9093]*kernel[3]+tmp[9094]*kernel[4]+tmp[9095]*kernel[5]+tmp[9193]*kernel[6]+tmp[9194]*kernel[7]+tmp[9195]*kernel[8];
				ans[9095]<=tmp[8994]*kernel[0]+tmp[8995]*kernel[1]+tmp[8996]*kernel[2]+tmp[9094]*kernel[3]+tmp[9095]*kernel[4]+tmp[9096]*kernel[5]+tmp[9194]*kernel[6]+tmp[9195]*kernel[7]+tmp[9196]*kernel[8];
				ans[9096]<=tmp[8995]*kernel[0]+tmp[8996]*kernel[1]+tmp[8997]*kernel[2]+tmp[9095]*kernel[3]+tmp[9096]*kernel[4]+tmp[9097]*kernel[5]+tmp[9195]*kernel[6]+tmp[9196]*kernel[7]+tmp[9197]*kernel[8];
				ans[9097]<=tmp[8996]*kernel[0]+tmp[8997]*kernel[1]+tmp[8998]*kernel[2]+tmp[9096]*kernel[3]+tmp[9097]*kernel[4]+tmp[9098]*kernel[5]+tmp[9196]*kernel[6]+tmp[9197]*kernel[7]+tmp[9198]*kernel[8];
				ans[9098]<=tmp[8997]*kernel[0]+tmp[8998]*kernel[1]+tmp[8999]*kernel[2]+tmp[9097]*kernel[3]+tmp[9098]*kernel[4]+tmp[9099]*kernel[5]+tmp[9197]*kernel[6]+tmp[9198]*kernel[7]+tmp[9199]*kernel[8];
				ans[9099]<=tmp[8998]*kernel[0]+tmp[8999]*kernel[1]+tmp[9098]*kernel[3]+tmp[9099]*kernel[4]+tmp[9198]*kernel[6]+tmp[9199]*kernel[7];
				ans[9100]<=tmp[9000]*kernel[1]+tmp[9001]*kernel[2]+tmp[9100]*kernel[4]+tmp[9101]*kernel[5]+tmp[9200]*kernel[7]+tmp[9201]*kernel[8];
				ans[9101]<=tmp[9000]*kernel[0]+tmp[9001]*kernel[1]+tmp[9002]*kernel[2]+tmp[9100]*kernel[3]+tmp[9101]*kernel[4]+tmp[9102]*kernel[5]+tmp[9200]*kernel[6]+tmp[9201]*kernel[7]+tmp[9202]*kernel[8];
				ans[9102]<=tmp[9001]*kernel[0]+tmp[9002]*kernel[1]+tmp[9003]*kernel[2]+tmp[9101]*kernel[3]+tmp[9102]*kernel[4]+tmp[9103]*kernel[5]+tmp[9201]*kernel[6]+tmp[9202]*kernel[7]+tmp[9203]*kernel[8];
				ans[9103]<=tmp[9002]*kernel[0]+tmp[9003]*kernel[1]+tmp[9004]*kernel[2]+tmp[9102]*kernel[3]+tmp[9103]*kernel[4]+tmp[9104]*kernel[5]+tmp[9202]*kernel[6]+tmp[9203]*kernel[7]+tmp[9204]*kernel[8];
				ans[9104]<=tmp[9003]*kernel[0]+tmp[9004]*kernel[1]+tmp[9005]*kernel[2]+tmp[9103]*kernel[3]+tmp[9104]*kernel[4]+tmp[9105]*kernel[5]+tmp[9203]*kernel[6]+tmp[9204]*kernel[7]+tmp[9205]*kernel[8];
				ans[9105]<=tmp[9004]*kernel[0]+tmp[9005]*kernel[1]+tmp[9006]*kernel[2]+tmp[9104]*kernel[3]+tmp[9105]*kernel[4]+tmp[9106]*kernel[5]+tmp[9204]*kernel[6]+tmp[9205]*kernel[7]+tmp[9206]*kernel[8];
				ans[9106]<=tmp[9005]*kernel[0]+tmp[9006]*kernel[1]+tmp[9007]*kernel[2]+tmp[9105]*kernel[3]+tmp[9106]*kernel[4]+tmp[9107]*kernel[5]+tmp[9205]*kernel[6]+tmp[9206]*kernel[7]+tmp[9207]*kernel[8];
				ans[9107]<=tmp[9006]*kernel[0]+tmp[9007]*kernel[1]+tmp[9008]*kernel[2]+tmp[9106]*kernel[3]+tmp[9107]*kernel[4]+tmp[9108]*kernel[5]+tmp[9206]*kernel[6]+tmp[9207]*kernel[7]+tmp[9208]*kernel[8];
				ans[9108]<=tmp[9007]*kernel[0]+tmp[9008]*kernel[1]+tmp[9009]*kernel[2]+tmp[9107]*kernel[3]+tmp[9108]*kernel[4]+tmp[9109]*kernel[5]+tmp[9207]*kernel[6]+tmp[9208]*kernel[7]+tmp[9209]*kernel[8];
				ans[9109]<=tmp[9008]*kernel[0]+tmp[9009]*kernel[1]+tmp[9010]*kernel[2]+tmp[9108]*kernel[3]+tmp[9109]*kernel[4]+tmp[9110]*kernel[5]+tmp[9208]*kernel[6]+tmp[9209]*kernel[7]+tmp[9210]*kernel[8];
				ans[9110]<=tmp[9009]*kernel[0]+tmp[9010]*kernel[1]+tmp[9011]*kernel[2]+tmp[9109]*kernel[3]+tmp[9110]*kernel[4]+tmp[9111]*kernel[5]+tmp[9209]*kernel[6]+tmp[9210]*kernel[7]+tmp[9211]*kernel[8];
				ans[9111]<=tmp[9010]*kernel[0]+tmp[9011]*kernel[1]+tmp[9012]*kernel[2]+tmp[9110]*kernel[3]+tmp[9111]*kernel[4]+tmp[9112]*kernel[5]+tmp[9210]*kernel[6]+tmp[9211]*kernel[7]+tmp[9212]*kernel[8];
				ans[9112]<=tmp[9011]*kernel[0]+tmp[9012]*kernel[1]+tmp[9013]*kernel[2]+tmp[9111]*kernel[3]+tmp[9112]*kernel[4]+tmp[9113]*kernel[5]+tmp[9211]*kernel[6]+tmp[9212]*kernel[7]+tmp[9213]*kernel[8];
				ans[9113]<=tmp[9012]*kernel[0]+tmp[9013]*kernel[1]+tmp[9014]*kernel[2]+tmp[9112]*kernel[3]+tmp[9113]*kernel[4]+tmp[9114]*kernel[5]+tmp[9212]*kernel[6]+tmp[9213]*kernel[7]+tmp[9214]*kernel[8];
				ans[9114]<=tmp[9013]*kernel[0]+tmp[9014]*kernel[1]+tmp[9015]*kernel[2]+tmp[9113]*kernel[3]+tmp[9114]*kernel[4]+tmp[9115]*kernel[5]+tmp[9213]*kernel[6]+tmp[9214]*kernel[7]+tmp[9215]*kernel[8];
				ans[9115]<=tmp[9014]*kernel[0]+tmp[9015]*kernel[1]+tmp[9016]*kernel[2]+tmp[9114]*kernel[3]+tmp[9115]*kernel[4]+tmp[9116]*kernel[5]+tmp[9214]*kernel[6]+tmp[9215]*kernel[7]+tmp[9216]*kernel[8];
				ans[9116]<=tmp[9015]*kernel[0]+tmp[9016]*kernel[1]+tmp[9017]*kernel[2]+tmp[9115]*kernel[3]+tmp[9116]*kernel[4]+tmp[9117]*kernel[5]+tmp[9215]*kernel[6]+tmp[9216]*kernel[7]+tmp[9217]*kernel[8];
				ans[9117]<=tmp[9016]*kernel[0]+tmp[9017]*kernel[1]+tmp[9018]*kernel[2]+tmp[9116]*kernel[3]+tmp[9117]*kernel[4]+tmp[9118]*kernel[5]+tmp[9216]*kernel[6]+tmp[9217]*kernel[7]+tmp[9218]*kernel[8];
				ans[9118]<=tmp[9017]*kernel[0]+tmp[9018]*kernel[1]+tmp[9019]*kernel[2]+tmp[9117]*kernel[3]+tmp[9118]*kernel[4]+tmp[9119]*kernel[5]+tmp[9217]*kernel[6]+tmp[9218]*kernel[7]+tmp[9219]*kernel[8];
				ans[9119]<=tmp[9018]*kernel[0]+tmp[9019]*kernel[1]+tmp[9020]*kernel[2]+tmp[9118]*kernel[3]+tmp[9119]*kernel[4]+tmp[9120]*kernel[5]+tmp[9218]*kernel[6]+tmp[9219]*kernel[7]+tmp[9220]*kernel[8];
				ans[9120]<=tmp[9019]*kernel[0]+tmp[9020]*kernel[1]+tmp[9021]*kernel[2]+tmp[9119]*kernel[3]+tmp[9120]*kernel[4]+tmp[9121]*kernel[5]+tmp[9219]*kernel[6]+tmp[9220]*kernel[7]+tmp[9221]*kernel[8];
				ans[9121]<=tmp[9020]*kernel[0]+tmp[9021]*kernel[1]+tmp[9022]*kernel[2]+tmp[9120]*kernel[3]+tmp[9121]*kernel[4]+tmp[9122]*kernel[5]+tmp[9220]*kernel[6]+tmp[9221]*kernel[7]+tmp[9222]*kernel[8];
				ans[9122]<=tmp[9021]*kernel[0]+tmp[9022]*kernel[1]+tmp[9023]*kernel[2]+tmp[9121]*kernel[3]+tmp[9122]*kernel[4]+tmp[9123]*kernel[5]+tmp[9221]*kernel[6]+tmp[9222]*kernel[7]+tmp[9223]*kernel[8];
				ans[9123]<=tmp[9022]*kernel[0]+tmp[9023]*kernel[1]+tmp[9024]*kernel[2]+tmp[9122]*kernel[3]+tmp[9123]*kernel[4]+tmp[9124]*kernel[5]+tmp[9222]*kernel[6]+tmp[9223]*kernel[7]+tmp[9224]*kernel[8];
				ans[9124]<=tmp[9023]*kernel[0]+tmp[9024]*kernel[1]+tmp[9025]*kernel[2]+tmp[9123]*kernel[3]+tmp[9124]*kernel[4]+tmp[9125]*kernel[5]+tmp[9223]*kernel[6]+tmp[9224]*kernel[7]+tmp[9225]*kernel[8];
				ans[9125]<=tmp[9024]*kernel[0]+tmp[9025]*kernel[1]+tmp[9026]*kernel[2]+tmp[9124]*kernel[3]+tmp[9125]*kernel[4]+tmp[9126]*kernel[5]+tmp[9224]*kernel[6]+tmp[9225]*kernel[7]+tmp[9226]*kernel[8];
				ans[9126]<=tmp[9025]*kernel[0]+tmp[9026]*kernel[1]+tmp[9027]*kernel[2]+tmp[9125]*kernel[3]+tmp[9126]*kernel[4]+tmp[9127]*kernel[5]+tmp[9225]*kernel[6]+tmp[9226]*kernel[7]+tmp[9227]*kernel[8];
				ans[9127]<=tmp[9026]*kernel[0]+tmp[9027]*kernel[1]+tmp[9028]*kernel[2]+tmp[9126]*kernel[3]+tmp[9127]*kernel[4]+tmp[9128]*kernel[5]+tmp[9226]*kernel[6]+tmp[9227]*kernel[7]+tmp[9228]*kernel[8];
				ans[9128]<=tmp[9027]*kernel[0]+tmp[9028]*kernel[1]+tmp[9029]*kernel[2]+tmp[9127]*kernel[3]+tmp[9128]*kernel[4]+tmp[9129]*kernel[5]+tmp[9227]*kernel[6]+tmp[9228]*kernel[7]+tmp[9229]*kernel[8];
				ans[9129]<=tmp[9028]*kernel[0]+tmp[9029]*kernel[1]+tmp[9030]*kernel[2]+tmp[9128]*kernel[3]+tmp[9129]*kernel[4]+tmp[9130]*kernel[5]+tmp[9228]*kernel[6]+tmp[9229]*kernel[7]+tmp[9230]*kernel[8];
				ans[9130]<=tmp[9029]*kernel[0]+tmp[9030]*kernel[1]+tmp[9031]*kernel[2]+tmp[9129]*kernel[3]+tmp[9130]*kernel[4]+tmp[9131]*kernel[5]+tmp[9229]*kernel[6]+tmp[9230]*kernel[7]+tmp[9231]*kernel[8];
				ans[9131]<=tmp[9030]*kernel[0]+tmp[9031]*kernel[1]+tmp[9032]*kernel[2]+tmp[9130]*kernel[3]+tmp[9131]*kernel[4]+tmp[9132]*kernel[5]+tmp[9230]*kernel[6]+tmp[9231]*kernel[7]+tmp[9232]*kernel[8];
				ans[9132]<=tmp[9031]*kernel[0]+tmp[9032]*kernel[1]+tmp[9033]*kernel[2]+tmp[9131]*kernel[3]+tmp[9132]*kernel[4]+tmp[9133]*kernel[5]+tmp[9231]*kernel[6]+tmp[9232]*kernel[7]+tmp[9233]*kernel[8];
				ans[9133]<=tmp[9032]*kernel[0]+tmp[9033]*kernel[1]+tmp[9034]*kernel[2]+tmp[9132]*kernel[3]+tmp[9133]*kernel[4]+tmp[9134]*kernel[5]+tmp[9232]*kernel[6]+tmp[9233]*kernel[7]+tmp[9234]*kernel[8];
				ans[9134]<=tmp[9033]*kernel[0]+tmp[9034]*kernel[1]+tmp[9035]*kernel[2]+tmp[9133]*kernel[3]+tmp[9134]*kernel[4]+tmp[9135]*kernel[5]+tmp[9233]*kernel[6]+tmp[9234]*kernel[7]+tmp[9235]*kernel[8];
				ans[9135]<=tmp[9034]*kernel[0]+tmp[9035]*kernel[1]+tmp[9036]*kernel[2]+tmp[9134]*kernel[3]+tmp[9135]*kernel[4]+tmp[9136]*kernel[5]+tmp[9234]*kernel[6]+tmp[9235]*kernel[7]+tmp[9236]*kernel[8];
				ans[9136]<=tmp[9035]*kernel[0]+tmp[9036]*kernel[1]+tmp[9037]*kernel[2]+tmp[9135]*kernel[3]+tmp[9136]*kernel[4]+tmp[9137]*kernel[5]+tmp[9235]*kernel[6]+tmp[9236]*kernel[7]+tmp[9237]*kernel[8];
				ans[9137]<=tmp[9036]*kernel[0]+tmp[9037]*kernel[1]+tmp[9038]*kernel[2]+tmp[9136]*kernel[3]+tmp[9137]*kernel[4]+tmp[9138]*kernel[5]+tmp[9236]*kernel[6]+tmp[9237]*kernel[7]+tmp[9238]*kernel[8];
				ans[9138]<=tmp[9037]*kernel[0]+tmp[9038]*kernel[1]+tmp[9039]*kernel[2]+tmp[9137]*kernel[3]+tmp[9138]*kernel[4]+tmp[9139]*kernel[5]+tmp[9237]*kernel[6]+tmp[9238]*kernel[7]+tmp[9239]*kernel[8];
				ans[9139]<=tmp[9038]*kernel[0]+tmp[9039]*kernel[1]+tmp[9040]*kernel[2]+tmp[9138]*kernel[3]+tmp[9139]*kernel[4]+tmp[9140]*kernel[5]+tmp[9238]*kernel[6]+tmp[9239]*kernel[7]+tmp[9240]*kernel[8];
				ans[9140]<=tmp[9039]*kernel[0]+tmp[9040]*kernel[1]+tmp[9041]*kernel[2]+tmp[9139]*kernel[3]+tmp[9140]*kernel[4]+tmp[9141]*kernel[5]+tmp[9239]*kernel[6]+tmp[9240]*kernel[7]+tmp[9241]*kernel[8];
				ans[9141]<=tmp[9040]*kernel[0]+tmp[9041]*kernel[1]+tmp[9042]*kernel[2]+tmp[9140]*kernel[3]+tmp[9141]*kernel[4]+tmp[9142]*kernel[5]+tmp[9240]*kernel[6]+tmp[9241]*kernel[7]+tmp[9242]*kernel[8];
				ans[9142]<=tmp[9041]*kernel[0]+tmp[9042]*kernel[1]+tmp[9043]*kernel[2]+tmp[9141]*kernel[3]+tmp[9142]*kernel[4]+tmp[9143]*kernel[5]+tmp[9241]*kernel[6]+tmp[9242]*kernel[7]+tmp[9243]*kernel[8];
				ans[9143]<=tmp[9042]*kernel[0]+tmp[9043]*kernel[1]+tmp[9044]*kernel[2]+tmp[9142]*kernel[3]+tmp[9143]*kernel[4]+tmp[9144]*kernel[5]+tmp[9242]*kernel[6]+tmp[9243]*kernel[7]+tmp[9244]*kernel[8];
				ans[9144]<=tmp[9043]*kernel[0]+tmp[9044]*kernel[1]+tmp[9045]*kernel[2]+tmp[9143]*kernel[3]+tmp[9144]*kernel[4]+tmp[9145]*kernel[5]+tmp[9243]*kernel[6]+tmp[9244]*kernel[7]+tmp[9245]*kernel[8];
				ans[9145]<=tmp[9044]*kernel[0]+tmp[9045]*kernel[1]+tmp[9046]*kernel[2]+tmp[9144]*kernel[3]+tmp[9145]*kernel[4]+tmp[9146]*kernel[5]+tmp[9244]*kernel[6]+tmp[9245]*kernel[7]+tmp[9246]*kernel[8];
				ans[9146]<=tmp[9045]*kernel[0]+tmp[9046]*kernel[1]+tmp[9047]*kernel[2]+tmp[9145]*kernel[3]+tmp[9146]*kernel[4]+tmp[9147]*kernel[5]+tmp[9245]*kernel[6]+tmp[9246]*kernel[7]+tmp[9247]*kernel[8];
				ans[9147]<=tmp[9046]*kernel[0]+tmp[9047]*kernel[1]+tmp[9048]*kernel[2]+tmp[9146]*kernel[3]+tmp[9147]*kernel[4]+tmp[9148]*kernel[5]+tmp[9246]*kernel[6]+tmp[9247]*kernel[7]+tmp[9248]*kernel[8];
				ans[9148]<=tmp[9047]*kernel[0]+tmp[9048]*kernel[1]+tmp[9049]*kernel[2]+tmp[9147]*kernel[3]+tmp[9148]*kernel[4]+tmp[9149]*kernel[5]+tmp[9247]*kernel[6]+tmp[9248]*kernel[7]+tmp[9249]*kernel[8];
				ans[9149]<=tmp[9048]*kernel[0]+tmp[9049]*kernel[1]+tmp[9050]*kernel[2]+tmp[9148]*kernel[3]+tmp[9149]*kernel[4]+tmp[9150]*kernel[5]+tmp[9248]*kernel[6]+tmp[9249]*kernel[7]+tmp[9250]*kernel[8];
				ans[9150]<=tmp[9049]*kernel[0]+tmp[9050]*kernel[1]+tmp[9051]*kernel[2]+tmp[9149]*kernel[3]+tmp[9150]*kernel[4]+tmp[9151]*kernel[5]+tmp[9249]*kernel[6]+tmp[9250]*kernel[7]+tmp[9251]*kernel[8];
				ans[9151]<=tmp[9050]*kernel[0]+tmp[9051]*kernel[1]+tmp[9052]*kernel[2]+tmp[9150]*kernel[3]+tmp[9151]*kernel[4]+tmp[9152]*kernel[5]+tmp[9250]*kernel[6]+tmp[9251]*kernel[7]+tmp[9252]*kernel[8];
				ans[9152]<=tmp[9051]*kernel[0]+tmp[9052]*kernel[1]+tmp[9053]*kernel[2]+tmp[9151]*kernel[3]+tmp[9152]*kernel[4]+tmp[9153]*kernel[5]+tmp[9251]*kernel[6]+tmp[9252]*kernel[7]+tmp[9253]*kernel[8];
				ans[9153]<=tmp[9052]*kernel[0]+tmp[9053]*kernel[1]+tmp[9054]*kernel[2]+tmp[9152]*kernel[3]+tmp[9153]*kernel[4]+tmp[9154]*kernel[5]+tmp[9252]*kernel[6]+tmp[9253]*kernel[7]+tmp[9254]*kernel[8];
				ans[9154]<=tmp[9053]*kernel[0]+tmp[9054]*kernel[1]+tmp[9055]*kernel[2]+tmp[9153]*kernel[3]+tmp[9154]*kernel[4]+tmp[9155]*kernel[5]+tmp[9253]*kernel[6]+tmp[9254]*kernel[7]+tmp[9255]*kernel[8];
				ans[9155]<=tmp[9054]*kernel[0]+tmp[9055]*kernel[1]+tmp[9056]*kernel[2]+tmp[9154]*kernel[3]+tmp[9155]*kernel[4]+tmp[9156]*kernel[5]+tmp[9254]*kernel[6]+tmp[9255]*kernel[7]+tmp[9256]*kernel[8];
				ans[9156]<=tmp[9055]*kernel[0]+tmp[9056]*kernel[1]+tmp[9057]*kernel[2]+tmp[9155]*kernel[3]+tmp[9156]*kernel[4]+tmp[9157]*kernel[5]+tmp[9255]*kernel[6]+tmp[9256]*kernel[7]+tmp[9257]*kernel[8];
				ans[9157]<=tmp[9056]*kernel[0]+tmp[9057]*kernel[1]+tmp[9058]*kernel[2]+tmp[9156]*kernel[3]+tmp[9157]*kernel[4]+tmp[9158]*kernel[5]+tmp[9256]*kernel[6]+tmp[9257]*kernel[7]+tmp[9258]*kernel[8];
				ans[9158]<=tmp[9057]*kernel[0]+tmp[9058]*kernel[1]+tmp[9059]*kernel[2]+tmp[9157]*kernel[3]+tmp[9158]*kernel[4]+tmp[9159]*kernel[5]+tmp[9257]*kernel[6]+tmp[9258]*kernel[7]+tmp[9259]*kernel[8];
				ans[9159]<=tmp[9058]*kernel[0]+tmp[9059]*kernel[1]+tmp[9060]*kernel[2]+tmp[9158]*kernel[3]+tmp[9159]*kernel[4]+tmp[9160]*kernel[5]+tmp[9258]*kernel[6]+tmp[9259]*kernel[7]+tmp[9260]*kernel[8];
				ans[9160]<=tmp[9059]*kernel[0]+tmp[9060]*kernel[1]+tmp[9061]*kernel[2]+tmp[9159]*kernel[3]+tmp[9160]*kernel[4]+tmp[9161]*kernel[5]+tmp[9259]*kernel[6]+tmp[9260]*kernel[7]+tmp[9261]*kernel[8];
				ans[9161]<=tmp[9060]*kernel[0]+tmp[9061]*kernel[1]+tmp[9062]*kernel[2]+tmp[9160]*kernel[3]+tmp[9161]*kernel[4]+tmp[9162]*kernel[5]+tmp[9260]*kernel[6]+tmp[9261]*kernel[7]+tmp[9262]*kernel[8];
				ans[9162]<=tmp[9061]*kernel[0]+tmp[9062]*kernel[1]+tmp[9063]*kernel[2]+tmp[9161]*kernel[3]+tmp[9162]*kernel[4]+tmp[9163]*kernel[5]+tmp[9261]*kernel[6]+tmp[9262]*kernel[7]+tmp[9263]*kernel[8];
				ans[9163]<=tmp[9062]*kernel[0]+tmp[9063]*kernel[1]+tmp[9064]*kernel[2]+tmp[9162]*kernel[3]+tmp[9163]*kernel[4]+tmp[9164]*kernel[5]+tmp[9262]*kernel[6]+tmp[9263]*kernel[7]+tmp[9264]*kernel[8];
				ans[9164]<=tmp[9063]*kernel[0]+tmp[9064]*kernel[1]+tmp[9065]*kernel[2]+tmp[9163]*kernel[3]+tmp[9164]*kernel[4]+tmp[9165]*kernel[5]+tmp[9263]*kernel[6]+tmp[9264]*kernel[7]+tmp[9265]*kernel[8];
				ans[9165]<=tmp[9064]*kernel[0]+tmp[9065]*kernel[1]+tmp[9066]*kernel[2]+tmp[9164]*kernel[3]+tmp[9165]*kernel[4]+tmp[9166]*kernel[5]+tmp[9264]*kernel[6]+tmp[9265]*kernel[7]+tmp[9266]*kernel[8];
				ans[9166]<=tmp[9065]*kernel[0]+tmp[9066]*kernel[1]+tmp[9067]*kernel[2]+tmp[9165]*kernel[3]+tmp[9166]*kernel[4]+tmp[9167]*kernel[5]+tmp[9265]*kernel[6]+tmp[9266]*kernel[7]+tmp[9267]*kernel[8];
				ans[9167]<=tmp[9066]*kernel[0]+tmp[9067]*kernel[1]+tmp[9068]*kernel[2]+tmp[9166]*kernel[3]+tmp[9167]*kernel[4]+tmp[9168]*kernel[5]+tmp[9266]*kernel[6]+tmp[9267]*kernel[7]+tmp[9268]*kernel[8];
				ans[9168]<=tmp[9067]*kernel[0]+tmp[9068]*kernel[1]+tmp[9069]*kernel[2]+tmp[9167]*kernel[3]+tmp[9168]*kernel[4]+tmp[9169]*kernel[5]+tmp[9267]*kernel[6]+tmp[9268]*kernel[7]+tmp[9269]*kernel[8];
				ans[9169]<=tmp[9068]*kernel[0]+tmp[9069]*kernel[1]+tmp[9070]*kernel[2]+tmp[9168]*kernel[3]+tmp[9169]*kernel[4]+tmp[9170]*kernel[5]+tmp[9268]*kernel[6]+tmp[9269]*kernel[7]+tmp[9270]*kernel[8];
				ans[9170]<=tmp[9069]*kernel[0]+tmp[9070]*kernel[1]+tmp[9071]*kernel[2]+tmp[9169]*kernel[3]+tmp[9170]*kernel[4]+tmp[9171]*kernel[5]+tmp[9269]*kernel[6]+tmp[9270]*kernel[7]+tmp[9271]*kernel[8];
				ans[9171]<=tmp[9070]*kernel[0]+tmp[9071]*kernel[1]+tmp[9072]*kernel[2]+tmp[9170]*kernel[3]+tmp[9171]*kernel[4]+tmp[9172]*kernel[5]+tmp[9270]*kernel[6]+tmp[9271]*kernel[7]+tmp[9272]*kernel[8];
				ans[9172]<=tmp[9071]*kernel[0]+tmp[9072]*kernel[1]+tmp[9073]*kernel[2]+tmp[9171]*kernel[3]+tmp[9172]*kernel[4]+tmp[9173]*kernel[5]+tmp[9271]*kernel[6]+tmp[9272]*kernel[7]+tmp[9273]*kernel[8];
				ans[9173]<=tmp[9072]*kernel[0]+tmp[9073]*kernel[1]+tmp[9074]*kernel[2]+tmp[9172]*kernel[3]+tmp[9173]*kernel[4]+tmp[9174]*kernel[5]+tmp[9272]*kernel[6]+tmp[9273]*kernel[7]+tmp[9274]*kernel[8];
				ans[9174]<=tmp[9073]*kernel[0]+tmp[9074]*kernel[1]+tmp[9075]*kernel[2]+tmp[9173]*kernel[3]+tmp[9174]*kernel[4]+tmp[9175]*kernel[5]+tmp[9273]*kernel[6]+tmp[9274]*kernel[7]+tmp[9275]*kernel[8];
				ans[9175]<=tmp[9074]*kernel[0]+tmp[9075]*kernel[1]+tmp[9076]*kernel[2]+tmp[9174]*kernel[3]+tmp[9175]*kernel[4]+tmp[9176]*kernel[5]+tmp[9274]*kernel[6]+tmp[9275]*kernel[7]+tmp[9276]*kernel[8];
				ans[9176]<=tmp[9075]*kernel[0]+tmp[9076]*kernel[1]+tmp[9077]*kernel[2]+tmp[9175]*kernel[3]+tmp[9176]*kernel[4]+tmp[9177]*kernel[5]+tmp[9275]*kernel[6]+tmp[9276]*kernel[7]+tmp[9277]*kernel[8];
				ans[9177]<=tmp[9076]*kernel[0]+tmp[9077]*kernel[1]+tmp[9078]*kernel[2]+tmp[9176]*kernel[3]+tmp[9177]*kernel[4]+tmp[9178]*kernel[5]+tmp[9276]*kernel[6]+tmp[9277]*kernel[7]+tmp[9278]*kernel[8];
				ans[9178]<=tmp[9077]*kernel[0]+tmp[9078]*kernel[1]+tmp[9079]*kernel[2]+tmp[9177]*kernel[3]+tmp[9178]*kernel[4]+tmp[9179]*kernel[5]+tmp[9277]*kernel[6]+tmp[9278]*kernel[7]+tmp[9279]*kernel[8];
				ans[9179]<=tmp[9078]*kernel[0]+tmp[9079]*kernel[1]+tmp[9080]*kernel[2]+tmp[9178]*kernel[3]+tmp[9179]*kernel[4]+tmp[9180]*kernel[5]+tmp[9278]*kernel[6]+tmp[9279]*kernel[7]+tmp[9280]*kernel[8];
				ans[9180]<=tmp[9079]*kernel[0]+tmp[9080]*kernel[1]+tmp[9081]*kernel[2]+tmp[9179]*kernel[3]+tmp[9180]*kernel[4]+tmp[9181]*kernel[5]+tmp[9279]*kernel[6]+tmp[9280]*kernel[7]+tmp[9281]*kernel[8];
				ans[9181]<=tmp[9080]*kernel[0]+tmp[9081]*kernel[1]+tmp[9082]*kernel[2]+tmp[9180]*kernel[3]+tmp[9181]*kernel[4]+tmp[9182]*kernel[5]+tmp[9280]*kernel[6]+tmp[9281]*kernel[7]+tmp[9282]*kernel[8];
				ans[9182]<=tmp[9081]*kernel[0]+tmp[9082]*kernel[1]+tmp[9083]*kernel[2]+tmp[9181]*kernel[3]+tmp[9182]*kernel[4]+tmp[9183]*kernel[5]+tmp[9281]*kernel[6]+tmp[9282]*kernel[7]+tmp[9283]*kernel[8];
				ans[9183]<=tmp[9082]*kernel[0]+tmp[9083]*kernel[1]+tmp[9084]*kernel[2]+tmp[9182]*kernel[3]+tmp[9183]*kernel[4]+tmp[9184]*kernel[5]+tmp[9282]*kernel[6]+tmp[9283]*kernel[7]+tmp[9284]*kernel[8];
				ans[9184]<=tmp[9083]*kernel[0]+tmp[9084]*kernel[1]+tmp[9085]*kernel[2]+tmp[9183]*kernel[3]+tmp[9184]*kernel[4]+tmp[9185]*kernel[5]+tmp[9283]*kernel[6]+tmp[9284]*kernel[7]+tmp[9285]*kernel[8];
				ans[9185]<=tmp[9084]*kernel[0]+tmp[9085]*kernel[1]+tmp[9086]*kernel[2]+tmp[9184]*kernel[3]+tmp[9185]*kernel[4]+tmp[9186]*kernel[5]+tmp[9284]*kernel[6]+tmp[9285]*kernel[7]+tmp[9286]*kernel[8];
				ans[9186]<=tmp[9085]*kernel[0]+tmp[9086]*kernel[1]+tmp[9087]*kernel[2]+tmp[9185]*kernel[3]+tmp[9186]*kernel[4]+tmp[9187]*kernel[5]+tmp[9285]*kernel[6]+tmp[9286]*kernel[7]+tmp[9287]*kernel[8];
				ans[9187]<=tmp[9086]*kernel[0]+tmp[9087]*kernel[1]+tmp[9088]*kernel[2]+tmp[9186]*kernel[3]+tmp[9187]*kernel[4]+tmp[9188]*kernel[5]+tmp[9286]*kernel[6]+tmp[9287]*kernel[7]+tmp[9288]*kernel[8];
				ans[9188]<=tmp[9087]*kernel[0]+tmp[9088]*kernel[1]+tmp[9089]*kernel[2]+tmp[9187]*kernel[3]+tmp[9188]*kernel[4]+tmp[9189]*kernel[5]+tmp[9287]*kernel[6]+tmp[9288]*kernel[7]+tmp[9289]*kernel[8];
				ans[9189]<=tmp[9088]*kernel[0]+tmp[9089]*kernel[1]+tmp[9090]*kernel[2]+tmp[9188]*kernel[3]+tmp[9189]*kernel[4]+tmp[9190]*kernel[5]+tmp[9288]*kernel[6]+tmp[9289]*kernel[7]+tmp[9290]*kernel[8];
				ans[9190]<=tmp[9089]*kernel[0]+tmp[9090]*kernel[1]+tmp[9091]*kernel[2]+tmp[9189]*kernel[3]+tmp[9190]*kernel[4]+tmp[9191]*kernel[5]+tmp[9289]*kernel[6]+tmp[9290]*kernel[7]+tmp[9291]*kernel[8];
				ans[9191]<=tmp[9090]*kernel[0]+tmp[9091]*kernel[1]+tmp[9092]*kernel[2]+tmp[9190]*kernel[3]+tmp[9191]*kernel[4]+tmp[9192]*kernel[5]+tmp[9290]*kernel[6]+tmp[9291]*kernel[7]+tmp[9292]*kernel[8];
				ans[9192]<=tmp[9091]*kernel[0]+tmp[9092]*kernel[1]+tmp[9093]*kernel[2]+tmp[9191]*kernel[3]+tmp[9192]*kernel[4]+tmp[9193]*kernel[5]+tmp[9291]*kernel[6]+tmp[9292]*kernel[7]+tmp[9293]*kernel[8];
				ans[9193]<=tmp[9092]*kernel[0]+tmp[9093]*kernel[1]+tmp[9094]*kernel[2]+tmp[9192]*kernel[3]+tmp[9193]*kernel[4]+tmp[9194]*kernel[5]+tmp[9292]*kernel[6]+tmp[9293]*kernel[7]+tmp[9294]*kernel[8];
				ans[9194]<=tmp[9093]*kernel[0]+tmp[9094]*kernel[1]+tmp[9095]*kernel[2]+tmp[9193]*kernel[3]+tmp[9194]*kernel[4]+tmp[9195]*kernel[5]+tmp[9293]*kernel[6]+tmp[9294]*kernel[7]+tmp[9295]*kernel[8];
				ans[9195]<=tmp[9094]*kernel[0]+tmp[9095]*kernel[1]+tmp[9096]*kernel[2]+tmp[9194]*kernel[3]+tmp[9195]*kernel[4]+tmp[9196]*kernel[5]+tmp[9294]*kernel[6]+tmp[9295]*kernel[7]+tmp[9296]*kernel[8];
				ans[9196]<=tmp[9095]*kernel[0]+tmp[9096]*kernel[1]+tmp[9097]*kernel[2]+tmp[9195]*kernel[3]+tmp[9196]*kernel[4]+tmp[9197]*kernel[5]+tmp[9295]*kernel[6]+tmp[9296]*kernel[7]+tmp[9297]*kernel[8];
				ans[9197]<=tmp[9096]*kernel[0]+tmp[9097]*kernel[1]+tmp[9098]*kernel[2]+tmp[9196]*kernel[3]+tmp[9197]*kernel[4]+tmp[9198]*kernel[5]+tmp[9296]*kernel[6]+tmp[9297]*kernel[7]+tmp[9298]*kernel[8];
				ans[9198]<=tmp[9097]*kernel[0]+tmp[9098]*kernel[1]+tmp[9099]*kernel[2]+tmp[9197]*kernel[3]+tmp[9198]*kernel[4]+tmp[9199]*kernel[5]+tmp[9297]*kernel[6]+tmp[9298]*kernel[7]+tmp[9299]*kernel[8];
				ans[9199]<=tmp[9098]*kernel[0]+tmp[9099]*kernel[1]+tmp[9198]*kernel[3]+tmp[9199]*kernel[4]+tmp[9298]*kernel[6]+tmp[9299]*kernel[7];
				ans[9200]<=tmp[9100]*kernel[1]+tmp[9101]*kernel[2]+tmp[9200]*kernel[4]+tmp[9201]*kernel[5]+tmp[9300]*kernel[7]+tmp[9301]*kernel[8];
				ans[9201]<=tmp[9100]*kernel[0]+tmp[9101]*kernel[1]+tmp[9102]*kernel[2]+tmp[9200]*kernel[3]+tmp[9201]*kernel[4]+tmp[9202]*kernel[5]+tmp[9300]*kernel[6]+tmp[9301]*kernel[7]+tmp[9302]*kernel[8];
				ans[9202]<=tmp[9101]*kernel[0]+tmp[9102]*kernel[1]+tmp[9103]*kernel[2]+tmp[9201]*kernel[3]+tmp[9202]*kernel[4]+tmp[9203]*kernel[5]+tmp[9301]*kernel[6]+tmp[9302]*kernel[7]+tmp[9303]*kernel[8];
				ans[9203]<=tmp[9102]*kernel[0]+tmp[9103]*kernel[1]+tmp[9104]*kernel[2]+tmp[9202]*kernel[3]+tmp[9203]*kernel[4]+tmp[9204]*kernel[5]+tmp[9302]*kernel[6]+tmp[9303]*kernel[7]+tmp[9304]*kernel[8];
				ans[9204]<=tmp[9103]*kernel[0]+tmp[9104]*kernel[1]+tmp[9105]*kernel[2]+tmp[9203]*kernel[3]+tmp[9204]*kernel[4]+tmp[9205]*kernel[5]+tmp[9303]*kernel[6]+tmp[9304]*kernel[7]+tmp[9305]*kernel[8];
				ans[9205]<=tmp[9104]*kernel[0]+tmp[9105]*kernel[1]+tmp[9106]*kernel[2]+tmp[9204]*kernel[3]+tmp[9205]*kernel[4]+tmp[9206]*kernel[5]+tmp[9304]*kernel[6]+tmp[9305]*kernel[7]+tmp[9306]*kernel[8];
				ans[9206]<=tmp[9105]*kernel[0]+tmp[9106]*kernel[1]+tmp[9107]*kernel[2]+tmp[9205]*kernel[3]+tmp[9206]*kernel[4]+tmp[9207]*kernel[5]+tmp[9305]*kernel[6]+tmp[9306]*kernel[7]+tmp[9307]*kernel[8];
				ans[9207]<=tmp[9106]*kernel[0]+tmp[9107]*kernel[1]+tmp[9108]*kernel[2]+tmp[9206]*kernel[3]+tmp[9207]*kernel[4]+tmp[9208]*kernel[5]+tmp[9306]*kernel[6]+tmp[9307]*kernel[7]+tmp[9308]*kernel[8];
				ans[9208]<=tmp[9107]*kernel[0]+tmp[9108]*kernel[1]+tmp[9109]*kernel[2]+tmp[9207]*kernel[3]+tmp[9208]*kernel[4]+tmp[9209]*kernel[5]+tmp[9307]*kernel[6]+tmp[9308]*kernel[7]+tmp[9309]*kernel[8];
				ans[9209]<=tmp[9108]*kernel[0]+tmp[9109]*kernel[1]+tmp[9110]*kernel[2]+tmp[9208]*kernel[3]+tmp[9209]*kernel[4]+tmp[9210]*kernel[5]+tmp[9308]*kernel[6]+tmp[9309]*kernel[7]+tmp[9310]*kernel[8];
				ans[9210]<=tmp[9109]*kernel[0]+tmp[9110]*kernel[1]+tmp[9111]*kernel[2]+tmp[9209]*kernel[3]+tmp[9210]*kernel[4]+tmp[9211]*kernel[5]+tmp[9309]*kernel[6]+tmp[9310]*kernel[7]+tmp[9311]*kernel[8];
				ans[9211]<=tmp[9110]*kernel[0]+tmp[9111]*kernel[1]+tmp[9112]*kernel[2]+tmp[9210]*kernel[3]+tmp[9211]*kernel[4]+tmp[9212]*kernel[5]+tmp[9310]*kernel[6]+tmp[9311]*kernel[7]+tmp[9312]*kernel[8];
				ans[9212]<=tmp[9111]*kernel[0]+tmp[9112]*kernel[1]+tmp[9113]*kernel[2]+tmp[9211]*kernel[3]+tmp[9212]*kernel[4]+tmp[9213]*kernel[5]+tmp[9311]*kernel[6]+tmp[9312]*kernel[7]+tmp[9313]*kernel[8];
				ans[9213]<=tmp[9112]*kernel[0]+tmp[9113]*kernel[1]+tmp[9114]*kernel[2]+tmp[9212]*kernel[3]+tmp[9213]*kernel[4]+tmp[9214]*kernel[5]+tmp[9312]*kernel[6]+tmp[9313]*kernel[7]+tmp[9314]*kernel[8];
				ans[9214]<=tmp[9113]*kernel[0]+tmp[9114]*kernel[1]+tmp[9115]*kernel[2]+tmp[9213]*kernel[3]+tmp[9214]*kernel[4]+tmp[9215]*kernel[5]+tmp[9313]*kernel[6]+tmp[9314]*kernel[7]+tmp[9315]*kernel[8];
				ans[9215]<=tmp[9114]*kernel[0]+tmp[9115]*kernel[1]+tmp[9116]*kernel[2]+tmp[9214]*kernel[3]+tmp[9215]*kernel[4]+tmp[9216]*kernel[5]+tmp[9314]*kernel[6]+tmp[9315]*kernel[7]+tmp[9316]*kernel[8];
				ans[9216]<=tmp[9115]*kernel[0]+tmp[9116]*kernel[1]+tmp[9117]*kernel[2]+tmp[9215]*kernel[3]+tmp[9216]*kernel[4]+tmp[9217]*kernel[5]+tmp[9315]*kernel[6]+tmp[9316]*kernel[7]+tmp[9317]*kernel[8];
				ans[9217]<=tmp[9116]*kernel[0]+tmp[9117]*kernel[1]+tmp[9118]*kernel[2]+tmp[9216]*kernel[3]+tmp[9217]*kernel[4]+tmp[9218]*kernel[5]+tmp[9316]*kernel[6]+tmp[9317]*kernel[7]+tmp[9318]*kernel[8];
				ans[9218]<=tmp[9117]*kernel[0]+tmp[9118]*kernel[1]+tmp[9119]*kernel[2]+tmp[9217]*kernel[3]+tmp[9218]*kernel[4]+tmp[9219]*kernel[5]+tmp[9317]*kernel[6]+tmp[9318]*kernel[7]+tmp[9319]*kernel[8];
				ans[9219]<=tmp[9118]*kernel[0]+tmp[9119]*kernel[1]+tmp[9120]*kernel[2]+tmp[9218]*kernel[3]+tmp[9219]*kernel[4]+tmp[9220]*kernel[5]+tmp[9318]*kernel[6]+tmp[9319]*kernel[7]+tmp[9320]*kernel[8];
				ans[9220]<=tmp[9119]*kernel[0]+tmp[9120]*kernel[1]+tmp[9121]*kernel[2]+tmp[9219]*kernel[3]+tmp[9220]*kernel[4]+tmp[9221]*kernel[5]+tmp[9319]*kernel[6]+tmp[9320]*kernel[7]+tmp[9321]*kernel[8];
				ans[9221]<=tmp[9120]*kernel[0]+tmp[9121]*kernel[1]+tmp[9122]*kernel[2]+tmp[9220]*kernel[3]+tmp[9221]*kernel[4]+tmp[9222]*kernel[5]+tmp[9320]*kernel[6]+tmp[9321]*kernel[7]+tmp[9322]*kernel[8];
				ans[9222]<=tmp[9121]*kernel[0]+tmp[9122]*kernel[1]+tmp[9123]*kernel[2]+tmp[9221]*kernel[3]+tmp[9222]*kernel[4]+tmp[9223]*kernel[5]+tmp[9321]*kernel[6]+tmp[9322]*kernel[7]+tmp[9323]*kernel[8];
				ans[9223]<=tmp[9122]*kernel[0]+tmp[9123]*kernel[1]+tmp[9124]*kernel[2]+tmp[9222]*kernel[3]+tmp[9223]*kernel[4]+tmp[9224]*kernel[5]+tmp[9322]*kernel[6]+tmp[9323]*kernel[7]+tmp[9324]*kernel[8];
				ans[9224]<=tmp[9123]*kernel[0]+tmp[9124]*kernel[1]+tmp[9125]*kernel[2]+tmp[9223]*kernel[3]+tmp[9224]*kernel[4]+tmp[9225]*kernel[5]+tmp[9323]*kernel[6]+tmp[9324]*kernel[7]+tmp[9325]*kernel[8];
				ans[9225]<=tmp[9124]*kernel[0]+tmp[9125]*kernel[1]+tmp[9126]*kernel[2]+tmp[9224]*kernel[3]+tmp[9225]*kernel[4]+tmp[9226]*kernel[5]+tmp[9324]*kernel[6]+tmp[9325]*kernel[7]+tmp[9326]*kernel[8];
				ans[9226]<=tmp[9125]*kernel[0]+tmp[9126]*kernel[1]+tmp[9127]*kernel[2]+tmp[9225]*kernel[3]+tmp[9226]*kernel[4]+tmp[9227]*kernel[5]+tmp[9325]*kernel[6]+tmp[9326]*kernel[7]+tmp[9327]*kernel[8];
				ans[9227]<=tmp[9126]*kernel[0]+tmp[9127]*kernel[1]+tmp[9128]*kernel[2]+tmp[9226]*kernel[3]+tmp[9227]*kernel[4]+tmp[9228]*kernel[5]+tmp[9326]*kernel[6]+tmp[9327]*kernel[7]+tmp[9328]*kernel[8];
				ans[9228]<=tmp[9127]*kernel[0]+tmp[9128]*kernel[1]+tmp[9129]*kernel[2]+tmp[9227]*kernel[3]+tmp[9228]*kernel[4]+tmp[9229]*kernel[5]+tmp[9327]*kernel[6]+tmp[9328]*kernel[7]+tmp[9329]*kernel[8];
				ans[9229]<=tmp[9128]*kernel[0]+tmp[9129]*kernel[1]+tmp[9130]*kernel[2]+tmp[9228]*kernel[3]+tmp[9229]*kernel[4]+tmp[9230]*kernel[5]+tmp[9328]*kernel[6]+tmp[9329]*kernel[7]+tmp[9330]*kernel[8];
				ans[9230]<=tmp[9129]*kernel[0]+tmp[9130]*kernel[1]+tmp[9131]*kernel[2]+tmp[9229]*kernel[3]+tmp[9230]*kernel[4]+tmp[9231]*kernel[5]+tmp[9329]*kernel[6]+tmp[9330]*kernel[7]+tmp[9331]*kernel[8];
				ans[9231]<=tmp[9130]*kernel[0]+tmp[9131]*kernel[1]+tmp[9132]*kernel[2]+tmp[9230]*kernel[3]+tmp[9231]*kernel[4]+tmp[9232]*kernel[5]+tmp[9330]*kernel[6]+tmp[9331]*kernel[7]+tmp[9332]*kernel[8];
				ans[9232]<=tmp[9131]*kernel[0]+tmp[9132]*kernel[1]+tmp[9133]*kernel[2]+tmp[9231]*kernel[3]+tmp[9232]*kernel[4]+tmp[9233]*kernel[5]+tmp[9331]*kernel[6]+tmp[9332]*kernel[7]+tmp[9333]*kernel[8];
				ans[9233]<=tmp[9132]*kernel[0]+tmp[9133]*kernel[1]+tmp[9134]*kernel[2]+tmp[9232]*kernel[3]+tmp[9233]*kernel[4]+tmp[9234]*kernel[5]+tmp[9332]*kernel[6]+tmp[9333]*kernel[7]+tmp[9334]*kernel[8];
				ans[9234]<=tmp[9133]*kernel[0]+tmp[9134]*kernel[1]+tmp[9135]*kernel[2]+tmp[9233]*kernel[3]+tmp[9234]*kernel[4]+tmp[9235]*kernel[5]+tmp[9333]*kernel[6]+tmp[9334]*kernel[7]+tmp[9335]*kernel[8];
				ans[9235]<=tmp[9134]*kernel[0]+tmp[9135]*kernel[1]+tmp[9136]*kernel[2]+tmp[9234]*kernel[3]+tmp[9235]*kernel[4]+tmp[9236]*kernel[5]+tmp[9334]*kernel[6]+tmp[9335]*kernel[7]+tmp[9336]*kernel[8];
				ans[9236]<=tmp[9135]*kernel[0]+tmp[9136]*kernel[1]+tmp[9137]*kernel[2]+tmp[9235]*kernel[3]+tmp[9236]*kernel[4]+tmp[9237]*kernel[5]+tmp[9335]*kernel[6]+tmp[9336]*kernel[7]+tmp[9337]*kernel[8];
				ans[9237]<=tmp[9136]*kernel[0]+tmp[9137]*kernel[1]+tmp[9138]*kernel[2]+tmp[9236]*kernel[3]+tmp[9237]*kernel[4]+tmp[9238]*kernel[5]+tmp[9336]*kernel[6]+tmp[9337]*kernel[7]+tmp[9338]*kernel[8];
				ans[9238]<=tmp[9137]*kernel[0]+tmp[9138]*kernel[1]+tmp[9139]*kernel[2]+tmp[9237]*kernel[3]+tmp[9238]*kernel[4]+tmp[9239]*kernel[5]+tmp[9337]*kernel[6]+tmp[9338]*kernel[7]+tmp[9339]*kernel[8];
				ans[9239]<=tmp[9138]*kernel[0]+tmp[9139]*kernel[1]+tmp[9140]*kernel[2]+tmp[9238]*kernel[3]+tmp[9239]*kernel[4]+tmp[9240]*kernel[5]+tmp[9338]*kernel[6]+tmp[9339]*kernel[7]+tmp[9340]*kernel[8];
				ans[9240]<=tmp[9139]*kernel[0]+tmp[9140]*kernel[1]+tmp[9141]*kernel[2]+tmp[9239]*kernel[3]+tmp[9240]*kernel[4]+tmp[9241]*kernel[5]+tmp[9339]*kernel[6]+tmp[9340]*kernel[7]+tmp[9341]*kernel[8];
				ans[9241]<=tmp[9140]*kernel[0]+tmp[9141]*kernel[1]+tmp[9142]*kernel[2]+tmp[9240]*kernel[3]+tmp[9241]*kernel[4]+tmp[9242]*kernel[5]+tmp[9340]*kernel[6]+tmp[9341]*kernel[7]+tmp[9342]*kernel[8];
				ans[9242]<=tmp[9141]*kernel[0]+tmp[9142]*kernel[1]+tmp[9143]*kernel[2]+tmp[9241]*kernel[3]+tmp[9242]*kernel[4]+tmp[9243]*kernel[5]+tmp[9341]*kernel[6]+tmp[9342]*kernel[7]+tmp[9343]*kernel[8];
				ans[9243]<=tmp[9142]*kernel[0]+tmp[9143]*kernel[1]+tmp[9144]*kernel[2]+tmp[9242]*kernel[3]+tmp[9243]*kernel[4]+tmp[9244]*kernel[5]+tmp[9342]*kernel[6]+tmp[9343]*kernel[7]+tmp[9344]*kernel[8];
				ans[9244]<=tmp[9143]*kernel[0]+tmp[9144]*kernel[1]+tmp[9145]*kernel[2]+tmp[9243]*kernel[3]+tmp[9244]*kernel[4]+tmp[9245]*kernel[5]+tmp[9343]*kernel[6]+tmp[9344]*kernel[7]+tmp[9345]*kernel[8];
				ans[9245]<=tmp[9144]*kernel[0]+tmp[9145]*kernel[1]+tmp[9146]*kernel[2]+tmp[9244]*kernel[3]+tmp[9245]*kernel[4]+tmp[9246]*kernel[5]+tmp[9344]*kernel[6]+tmp[9345]*kernel[7]+tmp[9346]*kernel[8];
				ans[9246]<=tmp[9145]*kernel[0]+tmp[9146]*kernel[1]+tmp[9147]*kernel[2]+tmp[9245]*kernel[3]+tmp[9246]*kernel[4]+tmp[9247]*kernel[5]+tmp[9345]*kernel[6]+tmp[9346]*kernel[7]+tmp[9347]*kernel[8];
				ans[9247]<=tmp[9146]*kernel[0]+tmp[9147]*kernel[1]+tmp[9148]*kernel[2]+tmp[9246]*kernel[3]+tmp[9247]*kernel[4]+tmp[9248]*kernel[5]+tmp[9346]*kernel[6]+tmp[9347]*kernel[7]+tmp[9348]*kernel[8];
				ans[9248]<=tmp[9147]*kernel[0]+tmp[9148]*kernel[1]+tmp[9149]*kernel[2]+tmp[9247]*kernel[3]+tmp[9248]*kernel[4]+tmp[9249]*kernel[5]+tmp[9347]*kernel[6]+tmp[9348]*kernel[7]+tmp[9349]*kernel[8];
				ans[9249]<=tmp[9148]*kernel[0]+tmp[9149]*kernel[1]+tmp[9150]*kernel[2]+tmp[9248]*kernel[3]+tmp[9249]*kernel[4]+tmp[9250]*kernel[5]+tmp[9348]*kernel[6]+tmp[9349]*kernel[7]+tmp[9350]*kernel[8];
				ans[9250]<=tmp[9149]*kernel[0]+tmp[9150]*kernel[1]+tmp[9151]*kernel[2]+tmp[9249]*kernel[3]+tmp[9250]*kernel[4]+tmp[9251]*kernel[5]+tmp[9349]*kernel[6]+tmp[9350]*kernel[7]+tmp[9351]*kernel[8];
				ans[9251]<=tmp[9150]*kernel[0]+tmp[9151]*kernel[1]+tmp[9152]*kernel[2]+tmp[9250]*kernel[3]+tmp[9251]*kernel[4]+tmp[9252]*kernel[5]+tmp[9350]*kernel[6]+tmp[9351]*kernel[7]+tmp[9352]*kernel[8];
				ans[9252]<=tmp[9151]*kernel[0]+tmp[9152]*kernel[1]+tmp[9153]*kernel[2]+tmp[9251]*kernel[3]+tmp[9252]*kernel[4]+tmp[9253]*kernel[5]+tmp[9351]*kernel[6]+tmp[9352]*kernel[7]+tmp[9353]*kernel[8];
				ans[9253]<=tmp[9152]*kernel[0]+tmp[9153]*kernel[1]+tmp[9154]*kernel[2]+tmp[9252]*kernel[3]+tmp[9253]*kernel[4]+tmp[9254]*kernel[5]+tmp[9352]*kernel[6]+tmp[9353]*kernel[7]+tmp[9354]*kernel[8];
				ans[9254]<=tmp[9153]*kernel[0]+tmp[9154]*kernel[1]+tmp[9155]*kernel[2]+tmp[9253]*kernel[3]+tmp[9254]*kernel[4]+tmp[9255]*kernel[5]+tmp[9353]*kernel[6]+tmp[9354]*kernel[7]+tmp[9355]*kernel[8];
				ans[9255]<=tmp[9154]*kernel[0]+tmp[9155]*kernel[1]+tmp[9156]*kernel[2]+tmp[9254]*kernel[3]+tmp[9255]*kernel[4]+tmp[9256]*kernel[5]+tmp[9354]*kernel[6]+tmp[9355]*kernel[7]+tmp[9356]*kernel[8];
				ans[9256]<=tmp[9155]*kernel[0]+tmp[9156]*kernel[1]+tmp[9157]*kernel[2]+tmp[9255]*kernel[3]+tmp[9256]*kernel[4]+tmp[9257]*kernel[5]+tmp[9355]*kernel[6]+tmp[9356]*kernel[7]+tmp[9357]*kernel[8];
				ans[9257]<=tmp[9156]*kernel[0]+tmp[9157]*kernel[1]+tmp[9158]*kernel[2]+tmp[9256]*kernel[3]+tmp[9257]*kernel[4]+tmp[9258]*kernel[5]+tmp[9356]*kernel[6]+tmp[9357]*kernel[7]+tmp[9358]*kernel[8];
				ans[9258]<=tmp[9157]*kernel[0]+tmp[9158]*kernel[1]+tmp[9159]*kernel[2]+tmp[9257]*kernel[3]+tmp[9258]*kernel[4]+tmp[9259]*kernel[5]+tmp[9357]*kernel[6]+tmp[9358]*kernel[7]+tmp[9359]*kernel[8];
				ans[9259]<=tmp[9158]*kernel[0]+tmp[9159]*kernel[1]+tmp[9160]*kernel[2]+tmp[9258]*kernel[3]+tmp[9259]*kernel[4]+tmp[9260]*kernel[5]+tmp[9358]*kernel[6]+tmp[9359]*kernel[7]+tmp[9360]*kernel[8];
				ans[9260]<=tmp[9159]*kernel[0]+tmp[9160]*kernel[1]+tmp[9161]*kernel[2]+tmp[9259]*kernel[3]+tmp[9260]*kernel[4]+tmp[9261]*kernel[5]+tmp[9359]*kernel[6]+tmp[9360]*kernel[7]+tmp[9361]*kernel[8];
				ans[9261]<=tmp[9160]*kernel[0]+tmp[9161]*kernel[1]+tmp[9162]*kernel[2]+tmp[9260]*kernel[3]+tmp[9261]*kernel[4]+tmp[9262]*kernel[5]+tmp[9360]*kernel[6]+tmp[9361]*kernel[7]+tmp[9362]*kernel[8];
				ans[9262]<=tmp[9161]*kernel[0]+tmp[9162]*kernel[1]+tmp[9163]*kernel[2]+tmp[9261]*kernel[3]+tmp[9262]*kernel[4]+tmp[9263]*kernel[5]+tmp[9361]*kernel[6]+tmp[9362]*kernel[7]+tmp[9363]*kernel[8];
				ans[9263]<=tmp[9162]*kernel[0]+tmp[9163]*kernel[1]+tmp[9164]*kernel[2]+tmp[9262]*kernel[3]+tmp[9263]*kernel[4]+tmp[9264]*kernel[5]+tmp[9362]*kernel[6]+tmp[9363]*kernel[7]+tmp[9364]*kernel[8];
				ans[9264]<=tmp[9163]*kernel[0]+tmp[9164]*kernel[1]+tmp[9165]*kernel[2]+tmp[9263]*kernel[3]+tmp[9264]*kernel[4]+tmp[9265]*kernel[5]+tmp[9363]*kernel[6]+tmp[9364]*kernel[7]+tmp[9365]*kernel[8];
				ans[9265]<=tmp[9164]*kernel[0]+tmp[9165]*kernel[1]+tmp[9166]*kernel[2]+tmp[9264]*kernel[3]+tmp[9265]*kernel[4]+tmp[9266]*kernel[5]+tmp[9364]*kernel[6]+tmp[9365]*kernel[7]+tmp[9366]*kernel[8];
				ans[9266]<=tmp[9165]*kernel[0]+tmp[9166]*kernel[1]+tmp[9167]*kernel[2]+tmp[9265]*kernel[3]+tmp[9266]*kernel[4]+tmp[9267]*kernel[5]+tmp[9365]*kernel[6]+tmp[9366]*kernel[7]+tmp[9367]*kernel[8];
				ans[9267]<=tmp[9166]*kernel[0]+tmp[9167]*kernel[1]+tmp[9168]*kernel[2]+tmp[9266]*kernel[3]+tmp[9267]*kernel[4]+tmp[9268]*kernel[5]+tmp[9366]*kernel[6]+tmp[9367]*kernel[7]+tmp[9368]*kernel[8];
				ans[9268]<=tmp[9167]*kernel[0]+tmp[9168]*kernel[1]+tmp[9169]*kernel[2]+tmp[9267]*kernel[3]+tmp[9268]*kernel[4]+tmp[9269]*kernel[5]+tmp[9367]*kernel[6]+tmp[9368]*kernel[7]+tmp[9369]*kernel[8];
				ans[9269]<=tmp[9168]*kernel[0]+tmp[9169]*kernel[1]+tmp[9170]*kernel[2]+tmp[9268]*kernel[3]+tmp[9269]*kernel[4]+tmp[9270]*kernel[5]+tmp[9368]*kernel[6]+tmp[9369]*kernel[7]+tmp[9370]*kernel[8];
				ans[9270]<=tmp[9169]*kernel[0]+tmp[9170]*kernel[1]+tmp[9171]*kernel[2]+tmp[9269]*kernel[3]+tmp[9270]*kernel[4]+tmp[9271]*kernel[5]+tmp[9369]*kernel[6]+tmp[9370]*kernel[7]+tmp[9371]*kernel[8];
				ans[9271]<=tmp[9170]*kernel[0]+tmp[9171]*kernel[1]+tmp[9172]*kernel[2]+tmp[9270]*kernel[3]+tmp[9271]*kernel[4]+tmp[9272]*kernel[5]+tmp[9370]*kernel[6]+tmp[9371]*kernel[7]+tmp[9372]*kernel[8];
				ans[9272]<=tmp[9171]*kernel[0]+tmp[9172]*kernel[1]+tmp[9173]*kernel[2]+tmp[9271]*kernel[3]+tmp[9272]*kernel[4]+tmp[9273]*kernel[5]+tmp[9371]*kernel[6]+tmp[9372]*kernel[7]+tmp[9373]*kernel[8];
				ans[9273]<=tmp[9172]*kernel[0]+tmp[9173]*kernel[1]+tmp[9174]*kernel[2]+tmp[9272]*kernel[3]+tmp[9273]*kernel[4]+tmp[9274]*kernel[5]+tmp[9372]*kernel[6]+tmp[9373]*kernel[7]+tmp[9374]*kernel[8];
				ans[9274]<=tmp[9173]*kernel[0]+tmp[9174]*kernel[1]+tmp[9175]*kernel[2]+tmp[9273]*kernel[3]+tmp[9274]*kernel[4]+tmp[9275]*kernel[5]+tmp[9373]*kernel[6]+tmp[9374]*kernel[7]+tmp[9375]*kernel[8];
				ans[9275]<=tmp[9174]*kernel[0]+tmp[9175]*kernel[1]+tmp[9176]*kernel[2]+tmp[9274]*kernel[3]+tmp[9275]*kernel[4]+tmp[9276]*kernel[5]+tmp[9374]*kernel[6]+tmp[9375]*kernel[7]+tmp[9376]*kernel[8];
				ans[9276]<=tmp[9175]*kernel[0]+tmp[9176]*kernel[1]+tmp[9177]*kernel[2]+tmp[9275]*kernel[3]+tmp[9276]*kernel[4]+tmp[9277]*kernel[5]+tmp[9375]*kernel[6]+tmp[9376]*kernel[7]+tmp[9377]*kernel[8];
				ans[9277]<=tmp[9176]*kernel[0]+tmp[9177]*kernel[1]+tmp[9178]*kernel[2]+tmp[9276]*kernel[3]+tmp[9277]*kernel[4]+tmp[9278]*kernel[5]+tmp[9376]*kernel[6]+tmp[9377]*kernel[7]+tmp[9378]*kernel[8];
				ans[9278]<=tmp[9177]*kernel[0]+tmp[9178]*kernel[1]+tmp[9179]*kernel[2]+tmp[9277]*kernel[3]+tmp[9278]*kernel[4]+tmp[9279]*kernel[5]+tmp[9377]*kernel[6]+tmp[9378]*kernel[7]+tmp[9379]*kernel[8];
				ans[9279]<=tmp[9178]*kernel[0]+tmp[9179]*kernel[1]+tmp[9180]*kernel[2]+tmp[9278]*kernel[3]+tmp[9279]*kernel[4]+tmp[9280]*kernel[5]+tmp[9378]*kernel[6]+tmp[9379]*kernel[7]+tmp[9380]*kernel[8];
				ans[9280]<=tmp[9179]*kernel[0]+tmp[9180]*kernel[1]+tmp[9181]*kernel[2]+tmp[9279]*kernel[3]+tmp[9280]*kernel[4]+tmp[9281]*kernel[5]+tmp[9379]*kernel[6]+tmp[9380]*kernel[7]+tmp[9381]*kernel[8];
				ans[9281]<=tmp[9180]*kernel[0]+tmp[9181]*kernel[1]+tmp[9182]*kernel[2]+tmp[9280]*kernel[3]+tmp[9281]*kernel[4]+tmp[9282]*kernel[5]+tmp[9380]*kernel[6]+tmp[9381]*kernel[7]+tmp[9382]*kernel[8];
				ans[9282]<=tmp[9181]*kernel[0]+tmp[9182]*kernel[1]+tmp[9183]*kernel[2]+tmp[9281]*kernel[3]+tmp[9282]*kernel[4]+tmp[9283]*kernel[5]+tmp[9381]*kernel[6]+tmp[9382]*kernel[7]+tmp[9383]*kernel[8];
				ans[9283]<=tmp[9182]*kernel[0]+tmp[9183]*kernel[1]+tmp[9184]*kernel[2]+tmp[9282]*kernel[3]+tmp[9283]*kernel[4]+tmp[9284]*kernel[5]+tmp[9382]*kernel[6]+tmp[9383]*kernel[7]+tmp[9384]*kernel[8];
				ans[9284]<=tmp[9183]*kernel[0]+tmp[9184]*kernel[1]+tmp[9185]*kernel[2]+tmp[9283]*kernel[3]+tmp[9284]*kernel[4]+tmp[9285]*kernel[5]+tmp[9383]*kernel[6]+tmp[9384]*kernel[7]+tmp[9385]*kernel[8];
				ans[9285]<=tmp[9184]*kernel[0]+tmp[9185]*kernel[1]+tmp[9186]*kernel[2]+tmp[9284]*kernel[3]+tmp[9285]*kernel[4]+tmp[9286]*kernel[5]+tmp[9384]*kernel[6]+tmp[9385]*kernel[7]+tmp[9386]*kernel[8];
				ans[9286]<=tmp[9185]*kernel[0]+tmp[9186]*kernel[1]+tmp[9187]*kernel[2]+tmp[9285]*kernel[3]+tmp[9286]*kernel[4]+tmp[9287]*kernel[5]+tmp[9385]*kernel[6]+tmp[9386]*kernel[7]+tmp[9387]*kernel[8];
				ans[9287]<=tmp[9186]*kernel[0]+tmp[9187]*kernel[1]+tmp[9188]*kernel[2]+tmp[9286]*kernel[3]+tmp[9287]*kernel[4]+tmp[9288]*kernel[5]+tmp[9386]*kernel[6]+tmp[9387]*kernel[7]+tmp[9388]*kernel[8];
				ans[9288]<=tmp[9187]*kernel[0]+tmp[9188]*kernel[1]+tmp[9189]*kernel[2]+tmp[9287]*kernel[3]+tmp[9288]*kernel[4]+tmp[9289]*kernel[5]+tmp[9387]*kernel[6]+tmp[9388]*kernel[7]+tmp[9389]*kernel[8];
				ans[9289]<=tmp[9188]*kernel[0]+tmp[9189]*kernel[1]+tmp[9190]*kernel[2]+tmp[9288]*kernel[3]+tmp[9289]*kernel[4]+tmp[9290]*kernel[5]+tmp[9388]*kernel[6]+tmp[9389]*kernel[7]+tmp[9390]*kernel[8];
				ans[9290]<=tmp[9189]*kernel[0]+tmp[9190]*kernel[1]+tmp[9191]*kernel[2]+tmp[9289]*kernel[3]+tmp[9290]*kernel[4]+tmp[9291]*kernel[5]+tmp[9389]*kernel[6]+tmp[9390]*kernel[7]+tmp[9391]*kernel[8];
				ans[9291]<=tmp[9190]*kernel[0]+tmp[9191]*kernel[1]+tmp[9192]*kernel[2]+tmp[9290]*kernel[3]+tmp[9291]*kernel[4]+tmp[9292]*kernel[5]+tmp[9390]*kernel[6]+tmp[9391]*kernel[7]+tmp[9392]*kernel[8];
				ans[9292]<=tmp[9191]*kernel[0]+tmp[9192]*kernel[1]+tmp[9193]*kernel[2]+tmp[9291]*kernel[3]+tmp[9292]*kernel[4]+tmp[9293]*kernel[5]+tmp[9391]*kernel[6]+tmp[9392]*kernel[7]+tmp[9393]*kernel[8];
				ans[9293]<=tmp[9192]*kernel[0]+tmp[9193]*kernel[1]+tmp[9194]*kernel[2]+tmp[9292]*kernel[3]+tmp[9293]*kernel[4]+tmp[9294]*kernel[5]+tmp[9392]*kernel[6]+tmp[9393]*kernel[7]+tmp[9394]*kernel[8];
				ans[9294]<=tmp[9193]*kernel[0]+tmp[9194]*kernel[1]+tmp[9195]*kernel[2]+tmp[9293]*kernel[3]+tmp[9294]*kernel[4]+tmp[9295]*kernel[5]+tmp[9393]*kernel[6]+tmp[9394]*kernel[7]+tmp[9395]*kernel[8];
				ans[9295]<=tmp[9194]*kernel[0]+tmp[9195]*kernel[1]+tmp[9196]*kernel[2]+tmp[9294]*kernel[3]+tmp[9295]*kernel[4]+tmp[9296]*kernel[5]+tmp[9394]*kernel[6]+tmp[9395]*kernel[7]+tmp[9396]*kernel[8];
				ans[9296]<=tmp[9195]*kernel[0]+tmp[9196]*kernel[1]+tmp[9197]*kernel[2]+tmp[9295]*kernel[3]+tmp[9296]*kernel[4]+tmp[9297]*kernel[5]+tmp[9395]*kernel[6]+tmp[9396]*kernel[7]+tmp[9397]*kernel[8];
				ans[9297]<=tmp[9196]*kernel[0]+tmp[9197]*kernel[1]+tmp[9198]*kernel[2]+tmp[9296]*kernel[3]+tmp[9297]*kernel[4]+tmp[9298]*kernel[5]+tmp[9396]*kernel[6]+tmp[9397]*kernel[7]+tmp[9398]*kernel[8];
				ans[9298]<=tmp[9197]*kernel[0]+tmp[9198]*kernel[1]+tmp[9199]*kernel[2]+tmp[9297]*kernel[3]+tmp[9298]*kernel[4]+tmp[9299]*kernel[5]+tmp[9397]*kernel[6]+tmp[9398]*kernel[7]+tmp[9399]*kernel[8];
				ans[9299]<=tmp[9198]*kernel[0]+tmp[9199]*kernel[1]+tmp[9298]*kernel[3]+tmp[9299]*kernel[4]+tmp[9398]*kernel[6]+tmp[9399]*kernel[7];
				ans[9300]<=tmp[9200]*kernel[1]+tmp[9201]*kernel[2]+tmp[9300]*kernel[4]+tmp[9301]*kernel[5]+tmp[9400]*kernel[7]+tmp[9401]*kernel[8];
				ans[9301]<=tmp[9200]*kernel[0]+tmp[9201]*kernel[1]+tmp[9202]*kernel[2]+tmp[9300]*kernel[3]+tmp[9301]*kernel[4]+tmp[9302]*kernel[5]+tmp[9400]*kernel[6]+tmp[9401]*kernel[7]+tmp[9402]*kernel[8];
				ans[9302]<=tmp[9201]*kernel[0]+tmp[9202]*kernel[1]+tmp[9203]*kernel[2]+tmp[9301]*kernel[3]+tmp[9302]*kernel[4]+tmp[9303]*kernel[5]+tmp[9401]*kernel[6]+tmp[9402]*kernel[7]+tmp[9403]*kernel[8];
				ans[9303]<=tmp[9202]*kernel[0]+tmp[9203]*kernel[1]+tmp[9204]*kernel[2]+tmp[9302]*kernel[3]+tmp[9303]*kernel[4]+tmp[9304]*kernel[5]+tmp[9402]*kernel[6]+tmp[9403]*kernel[7]+tmp[9404]*kernel[8];
				ans[9304]<=tmp[9203]*kernel[0]+tmp[9204]*kernel[1]+tmp[9205]*kernel[2]+tmp[9303]*kernel[3]+tmp[9304]*kernel[4]+tmp[9305]*kernel[5]+tmp[9403]*kernel[6]+tmp[9404]*kernel[7]+tmp[9405]*kernel[8];
				ans[9305]<=tmp[9204]*kernel[0]+tmp[9205]*kernel[1]+tmp[9206]*kernel[2]+tmp[9304]*kernel[3]+tmp[9305]*kernel[4]+tmp[9306]*kernel[5]+tmp[9404]*kernel[6]+tmp[9405]*kernel[7]+tmp[9406]*kernel[8];
				ans[9306]<=tmp[9205]*kernel[0]+tmp[9206]*kernel[1]+tmp[9207]*kernel[2]+tmp[9305]*kernel[3]+tmp[9306]*kernel[4]+tmp[9307]*kernel[5]+tmp[9405]*kernel[6]+tmp[9406]*kernel[7]+tmp[9407]*kernel[8];
				ans[9307]<=tmp[9206]*kernel[0]+tmp[9207]*kernel[1]+tmp[9208]*kernel[2]+tmp[9306]*kernel[3]+tmp[9307]*kernel[4]+tmp[9308]*kernel[5]+tmp[9406]*kernel[6]+tmp[9407]*kernel[7]+tmp[9408]*kernel[8];
				ans[9308]<=tmp[9207]*kernel[0]+tmp[9208]*kernel[1]+tmp[9209]*kernel[2]+tmp[9307]*kernel[3]+tmp[9308]*kernel[4]+tmp[9309]*kernel[5]+tmp[9407]*kernel[6]+tmp[9408]*kernel[7]+tmp[9409]*kernel[8];
				ans[9309]<=tmp[9208]*kernel[0]+tmp[9209]*kernel[1]+tmp[9210]*kernel[2]+tmp[9308]*kernel[3]+tmp[9309]*kernel[4]+tmp[9310]*kernel[5]+tmp[9408]*kernel[6]+tmp[9409]*kernel[7]+tmp[9410]*kernel[8];
				ans[9310]<=tmp[9209]*kernel[0]+tmp[9210]*kernel[1]+tmp[9211]*kernel[2]+tmp[9309]*kernel[3]+tmp[9310]*kernel[4]+tmp[9311]*kernel[5]+tmp[9409]*kernel[6]+tmp[9410]*kernel[7]+tmp[9411]*kernel[8];
				ans[9311]<=tmp[9210]*kernel[0]+tmp[9211]*kernel[1]+tmp[9212]*kernel[2]+tmp[9310]*kernel[3]+tmp[9311]*kernel[4]+tmp[9312]*kernel[5]+tmp[9410]*kernel[6]+tmp[9411]*kernel[7]+tmp[9412]*kernel[8];
				ans[9312]<=tmp[9211]*kernel[0]+tmp[9212]*kernel[1]+tmp[9213]*kernel[2]+tmp[9311]*kernel[3]+tmp[9312]*kernel[4]+tmp[9313]*kernel[5]+tmp[9411]*kernel[6]+tmp[9412]*kernel[7]+tmp[9413]*kernel[8];
				ans[9313]<=tmp[9212]*kernel[0]+tmp[9213]*kernel[1]+tmp[9214]*kernel[2]+tmp[9312]*kernel[3]+tmp[9313]*kernel[4]+tmp[9314]*kernel[5]+tmp[9412]*kernel[6]+tmp[9413]*kernel[7]+tmp[9414]*kernel[8];
				ans[9314]<=tmp[9213]*kernel[0]+tmp[9214]*kernel[1]+tmp[9215]*kernel[2]+tmp[9313]*kernel[3]+tmp[9314]*kernel[4]+tmp[9315]*kernel[5]+tmp[9413]*kernel[6]+tmp[9414]*kernel[7]+tmp[9415]*kernel[8];
				ans[9315]<=tmp[9214]*kernel[0]+tmp[9215]*kernel[1]+tmp[9216]*kernel[2]+tmp[9314]*kernel[3]+tmp[9315]*kernel[4]+tmp[9316]*kernel[5]+tmp[9414]*kernel[6]+tmp[9415]*kernel[7]+tmp[9416]*kernel[8];
				ans[9316]<=tmp[9215]*kernel[0]+tmp[9216]*kernel[1]+tmp[9217]*kernel[2]+tmp[9315]*kernel[3]+tmp[9316]*kernel[4]+tmp[9317]*kernel[5]+tmp[9415]*kernel[6]+tmp[9416]*kernel[7]+tmp[9417]*kernel[8];
				ans[9317]<=tmp[9216]*kernel[0]+tmp[9217]*kernel[1]+tmp[9218]*kernel[2]+tmp[9316]*kernel[3]+tmp[9317]*kernel[4]+tmp[9318]*kernel[5]+tmp[9416]*kernel[6]+tmp[9417]*kernel[7]+tmp[9418]*kernel[8];
				ans[9318]<=tmp[9217]*kernel[0]+tmp[9218]*kernel[1]+tmp[9219]*kernel[2]+tmp[9317]*kernel[3]+tmp[9318]*kernel[4]+tmp[9319]*kernel[5]+tmp[9417]*kernel[6]+tmp[9418]*kernel[7]+tmp[9419]*kernel[8];
				ans[9319]<=tmp[9218]*kernel[0]+tmp[9219]*kernel[1]+tmp[9220]*kernel[2]+tmp[9318]*kernel[3]+tmp[9319]*kernel[4]+tmp[9320]*kernel[5]+tmp[9418]*kernel[6]+tmp[9419]*kernel[7]+tmp[9420]*kernel[8];
				ans[9320]<=tmp[9219]*kernel[0]+tmp[9220]*kernel[1]+tmp[9221]*kernel[2]+tmp[9319]*kernel[3]+tmp[9320]*kernel[4]+tmp[9321]*kernel[5]+tmp[9419]*kernel[6]+tmp[9420]*kernel[7]+tmp[9421]*kernel[8];
				ans[9321]<=tmp[9220]*kernel[0]+tmp[9221]*kernel[1]+tmp[9222]*kernel[2]+tmp[9320]*kernel[3]+tmp[9321]*kernel[4]+tmp[9322]*kernel[5]+tmp[9420]*kernel[6]+tmp[9421]*kernel[7]+tmp[9422]*kernel[8];
				ans[9322]<=tmp[9221]*kernel[0]+tmp[9222]*kernel[1]+tmp[9223]*kernel[2]+tmp[9321]*kernel[3]+tmp[9322]*kernel[4]+tmp[9323]*kernel[5]+tmp[9421]*kernel[6]+tmp[9422]*kernel[7]+tmp[9423]*kernel[8];
				ans[9323]<=tmp[9222]*kernel[0]+tmp[9223]*kernel[1]+tmp[9224]*kernel[2]+tmp[9322]*kernel[3]+tmp[9323]*kernel[4]+tmp[9324]*kernel[5]+tmp[9422]*kernel[6]+tmp[9423]*kernel[7]+tmp[9424]*kernel[8];
				ans[9324]<=tmp[9223]*kernel[0]+tmp[9224]*kernel[1]+tmp[9225]*kernel[2]+tmp[9323]*kernel[3]+tmp[9324]*kernel[4]+tmp[9325]*kernel[5]+tmp[9423]*kernel[6]+tmp[9424]*kernel[7]+tmp[9425]*kernel[8];
				ans[9325]<=tmp[9224]*kernel[0]+tmp[9225]*kernel[1]+tmp[9226]*kernel[2]+tmp[9324]*kernel[3]+tmp[9325]*kernel[4]+tmp[9326]*kernel[5]+tmp[9424]*kernel[6]+tmp[9425]*kernel[7]+tmp[9426]*kernel[8];
				ans[9326]<=tmp[9225]*kernel[0]+tmp[9226]*kernel[1]+tmp[9227]*kernel[2]+tmp[9325]*kernel[3]+tmp[9326]*kernel[4]+tmp[9327]*kernel[5]+tmp[9425]*kernel[6]+tmp[9426]*kernel[7]+tmp[9427]*kernel[8];
				ans[9327]<=tmp[9226]*kernel[0]+tmp[9227]*kernel[1]+tmp[9228]*kernel[2]+tmp[9326]*kernel[3]+tmp[9327]*kernel[4]+tmp[9328]*kernel[5]+tmp[9426]*kernel[6]+tmp[9427]*kernel[7]+tmp[9428]*kernel[8];
				ans[9328]<=tmp[9227]*kernel[0]+tmp[9228]*kernel[1]+tmp[9229]*kernel[2]+tmp[9327]*kernel[3]+tmp[9328]*kernel[4]+tmp[9329]*kernel[5]+tmp[9427]*kernel[6]+tmp[9428]*kernel[7]+tmp[9429]*kernel[8];
				ans[9329]<=tmp[9228]*kernel[0]+tmp[9229]*kernel[1]+tmp[9230]*kernel[2]+tmp[9328]*kernel[3]+tmp[9329]*kernel[4]+tmp[9330]*kernel[5]+tmp[9428]*kernel[6]+tmp[9429]*kernel[7]+tmp[9430]*kernel[8];
				ans[9330]<=tmp[9229]*kernel[0]+tmp[9230]*kernel[1]+tmp[9231]*kernel[2]+tmp[9329]*kernel[3]+tmp[9330]*kernel[4]+tmp[9331]*kernel[5]+tmp[9429]*kernel[6]+tmp[9430]*kernel[7]+tmp[9431]*kernel[8];
				ans[9331]<=tmp[9230]*kernel[0]+tmp[9231]*kernel[1]+tmp[9232]*kernel[2]+tmp[9330]*kernel[3]+tmp[9331]*kernel[4]+tmp[9332]*kernel[5]+tmp[9430]*kernel[6]+tmp[9431]*kernel[7]+tmp[9432]*kernel[8];
				ans[9332]<=tmp[9231]*kernel[0]+tmp[9232]*kernel[1]+tmp[9233]*kernel[2]+tmp[9331]*kernel[3]+tmp[9332]*kernel[4]+tmp[9333]*kernel[5]+tmp[9431]*kernel[6]+tmp[9432]*kernel[7]+tmp[9433]*kernel[8];
				ans[9333]<=tmp[9232]*kernel[0]+tmp[9233]*kernel[1]+tmp[9234]*kernel[2]+tmp[9332]*kernel[3]+tmp[9333]*kernel[4]+tmp[9334]*kernel[5]+tmp[9432]*kernel[6]+tmp[9433]*kernel[7]+tmp[9434]*kernel[8];
				ans[9334]<=tmp[9233]*kernel[0]+tmp[9234]*kernel[1]+tmp[9235]*kernel[2]+tmp[9333]*kernel[3]+tmp[9334]*kernel[4]+tmp[9335]*kernel[5]+tmp[9433]*kernel[6]+tmp[9434]*kernel[7]+tmp[9435]*kernel[8];
				ans[9335]<=tmp[9234]*kernel[0]+tmp[9235]*kernel[1]+tmp[9236]*kernel[2]+tmp[9334]*kernel[3]+tmp[9335]*kernel[4]+tmp[9336]*kernel[5]+tmp[9434]*kernel[6]+tmp[9435]*kernel[7]+tmp[9436]*kernel[8];
				ans[9336]<=tmp[9235]*kernel[0]+tmp[9236]*kernel[1]+tmp[9237]*kernel[2]+tmp[9335]*kernel[3]+tmp[9336]*kernel[4]+tmp[9337]*kernel[5]+tmp[9435]*kernel[6]+tmp[9436]*kernel[7]+tmp[9437]*kernel[8];
				ans[9337]<=tmp[9236]*kernel[0]+tmp[9237]*kernel[1]+tmp[9238]*kernel[2]+tmp[9336]*kernel[3]+tmp[9337]*kernel[4]+tmp[9338]*kernel[5]+tmp[9436]*kernel[6]+tmp[9437]*kernel[7]+tmp[9438]*kernel[8];
				ans[9338]<=tmp[9237]*kernel[0]+tmp[9238]*kernel[1]+tmp[9239]*kernel[2]+tmp[9337]*kernel[3]+tmp[9338]*kernel[4]+tmp[9339]*kernel[5]+tmp[9437]*kernel[6]+tmp[9438]*kernel[7]+tmp[9439]*kernel[8];
				ans[9339]<=tmp[9238]*kernel[0]+tmp[9239]*kernel[1]+tmp[9240]*kernel[2]+tmp[9338]*kernel[3]+tmp[9339]*kernel[4]+tmp[9340]*kernel[5]+tmp[9438]*kernel[6]+tmp[9439]*kernel[7]+tmp[9440]*kernel[8];
				ans[9340]<=tmp[9239]*kernel[0]+tmp[9240]*kernel[1]+tmp[9241]*kernel[2]+tmp[9339]*kernel[3]+tmp[9340]*kernel[4]+tmp[9341]*kernel[5]+tmp[9439]*kernel[6]+tmp[9440]*kernel[7]+tmp[9441]*kernel[8];
				ans[9341]<=tmp[9240]*kernel[0]+tmp[9241]*kernel[1]+tmp[9242]*kernel[2]+tmp[9340]*kernel[3]+tmp[9341]*kernel[4]+tmp[9342]*kernel[5]+tmp[9440]*kernel[6]+tmp[9441]*kernel[7]+tmp[9442]*kernel[8];
				ans[9342]<=tmp[9241]*kernel[0]+tmp[9242]*kernel[1]+tmp[9243]*kernel[2]+tmp[9341]*kernel[3]+tmp[9342]*kernel[4]+tmp[9343]*kernel[5]+tmp[9441]*kernel[6]+tmp[9442]*kernel[7]+tmp[9443]*kernel[8];
				ans[9343]<=tmp[9242]*kernel[0]+tmp[9243]*kernel[1]+tmp[9244]*kernel[2]+tmp[9342]*kernel[3]+tmp[9343]*kernel[4]+tmp[9344]*kernel[5]+tmp[9442]*kernel[6]+tmp[9443]*kernel[7]+tmp[9444]*kernel[8];
				ans[9344]<=tmp[9243]*kernel[0]+tmp[9244]*kernel[1]+tmp[9245]*kernel[2]+tmp[9343]*kernel[3]+tmp[9344]*kernel[4]+tmp[9345]*kernel[5]+tmp[9443]*kernel[6]+tmp[9444]*kernel[7]+tmp[9445]*kernel[8];
				ans[9345]<=tmp[9244]*kernel[0]+tmp[9245]*kernel[1]+tmp[9246]*kernel[2]+tmp[9344]*kernel[3]+tmp[9345]*kernel[4]+tmp[9346]*kernel[5]+tmp[9444]*kernel[6]+tmp[9445]*kernel[7]+tmp[9446]*kernel[8];
				ans[9346]<=tmp[9245]*kernel[0]+tmp[9246]*kernel[1]+tmp[9247]*kernel[2]+tmp[9345]*kernel[3]+tmp[9346]*kernel[4]+tmp[9347]*kernel[5]+tmp[9445]*kernel[6]+tmp[9446]*kernel[7]+tmp[9447]*kernel[8];
				ans[9347]<=tmp[9246]*kernel[0]+tmp[9247]*kernel[1]+tmp[9248]*kernel[2]+tmp[9346]*kernel[3]+tmp[9347]*kernel[4]+tmp[9348]*kernel[5]+tmp[9446]*kernel[6]+tmp[9447]*kernel[7]+tmp[9448]*kernel[8];
				ans[9348]<=tmp[9247]*kernel[0]+tmp[9248]*kernel[1]+tmp[9249]*kernel[2]+tmp[9347]*kernel[3]+tmp[9348]*kernel[4]+tmp[9349]*kernel[5]+tmp[9447]*kernel[6]+tmp[9448]*kernel[7]+tmp[9449]*kernel[8];
				ans[9349]<=tmp[9248]*kernel[0]+tmp[9249]*kernel[1]+tmp[9250]*kernel[2]+tmp[9348]*kernel[3]+tmp[9349]*kernel[4]+tmp[9350]*kernel[5]+tmp[9448]*kernel[6]+tmp[9449]*kernel[7]+tmp[9450]*kernel[8];
				ans[9350]<=tmp[9249]*kernel[0]+tmp[9250]*kernel[1]+tmp[9251]*kernel[2]+tmp[9349]*kernel[3]+tmp[9350]*kernel[4]+tmp[9351]*kernel[5]+tmp[9449]*kernel[6]+tmp[9450]*kernel[7]+tmp[9451]*kernel[8];
				ans[9351]<=tmp[9250]*kernel[0]+tmp[9251]*kernel[1]+tmp[9252]*kernel[2]+tmp[9350]*kernel[3]+tmp[9351]*kernel[4]+tmp[9352]*kernel[5]+tmp[9450]*kernel[6]+tmp[9451]*kernel[7]+tmp[9452]*kernel[8];
				ans[9352]<=tmp[9251]*kernel[0]+tmp[9252]*kernel[1]+tmp[9253]*kernel[2]+tmp[9351]*kernel[3]+tmp[9352]*kernel[4]+tmp[9353]*kernel[5]+tmp[9451]*kernel[6]+tmp[9452]*kernel[7]+tmp[9453]*kernel[8];
				ans[9353]<=tmp[9252]*kernel[0]+tmp[9253]*kernel[1]+tmp[9254]*kernel[2]+tmp[9352]*kernel[3]+tmp[9353]*kernel[4]+tmp[9354]*kernel[5]+tmp[9452]*kernel[6]+tmp[9453]*kernel[7]+tmp[9454]*kernel[8];
				ans[9354]<=tmp[9253]*kernel[0]+tmp[9254]*kernel[1]+tmp[9255]*kernel[2]+tmp[9353]*kernel[3]+tmp[9354]*kernel[4]+tmp[9355]*kernel[5]+tmp[9453]*kernel[6]+tmp[9454]*kernel[7]+tmp[9455]*kernel[8];
				ans[9355]<=tmp[9254]*kernel[0]+tmp[9255]*kernel[1]+tmp[9256]*kernel[2]+tmp[9354]*kernel[3]+tmp[9355]*kernel[4]+tmp[9356]*kernel[5]+tmp[9454]*kernel[6]+tmp[9455]*kernel[7]+tmp[9456]*kernel[8];
				ans[9356]<=tmp[9255]*kernel[0]+tmp[9256]*kernel[1]+tmp[9257]*kernel[2]+tmp[9355]*kernel[3]+tmp[9356]*kernel[4]+tmp[9357]*kernel[5]+tmp[9455]*kernel[6]+tmp[9456]*kernel[7]+tmp[9457]*kernel[8];
				ans[9357]<=tmp[9256]*kernel[0]+tmp[9257]*kernel[1]+tmp[9258]*kernel[2]+tmp[9356]*kernel[3]+tmp[9357]*kernel[4]+tmp[9358]*kernel[5]+tmp[9456]*kernel[6]+tmp[9457]*kernel[7]+tmp[9458]*kernel[8];
				ans[9358]<=tmp[9257]*kernel[0]+tmp[9258]*kernel[1]+tmp[9259]*kernel[2]+tmp[9357]*kernel[3]+tmp[9358]*kernel[4]+tmp[9359]*kernel[5]+tmp[9457]*kernel[6]+tmp[9458]*kernel[7]+tmp[9459]*kernel[8];
				ans[9359]<=tmp[9258]*kernel[0]+tmp[9259]*kernel[1]+tmp[9260]*kernel[2]+tmp[9358]*kernel[3]+tmp[9359]*kernel[4]+tmp[9360]*kernel[5]+tmp[9458]*kernel[6]+tmp[9459]*kernel[7]+tmp[9460]*kernel[8];
				ans[9360]<=tmp[9259]*kernel[0]+tmp[9260]*kernel[1]+tmp[9261]*kernel[2]+tmp[9359]*kernel[3]+tmp[9360]*kernel[4]+tmp[9361]*kernel[5]+tmp[9459]*kernel[6]+tmp[9460]*kernel[7]+tmp[9461]*kernel[8];
				ans[9361]<=tmp[9260]*kernel[0]+tmp[9261]*kernel[1]+tmp[9262]*kernel[2]+tmp[9360]*kernel[3]+tmp[9361]*kernel[4]+tmp[9362]*kernel[5]+tmp[9460]*kernel[6]+tmp[9461]*kernel[7]+tmp[9462]*kernel[8];
				ans[9362]<=tmp[9261]*kernel[0]+tmp[9262]*kernel[1]+tmp[9263]*kernel[2]+tmp[9361]*kernel[3]+tmp[9362]*kernel[4]+tmp[9363]*kernel[5]+tmp[9461]*kernel[6]+tmp[9462]*kernel[7]+tmp[9463]*kernel[8];
				ans[9363]<=tmp[9262]*kernel[0]+tmp[9263]*kernel[1]+tmp[9264]*kernel[2]+tmp[9362]*kernel[3]+tmp[9363]*kernel[4]+tmp[9364]*kernel[5]+tmp[9462]*kernel[6]+tmp[9463]*kernel[7]+tmp[9464]*kernel[8];
				ans[9364]<=tmp[9263]*kernel[0]+tmp[9264]*kernel[1]+tmp[9265]*kernel[2]+tmp[9363]*kernel[3]+tmp[9364]*kernel[4]+tmp[9365]*kernel[5]+tmp[9463]*kernel[6]+tmp[9464]*kernel[7]+tmp[9465]*kernel[8];
				ans[9365]<=tmp[9264]*kernel[0]+tmp[9265]*kernel[1]+tmp[9266]*kernel[2]+tmp[9364]*kernel[3]+tmp[9365]*kernel[4]+tmp[9366]*kernel[5]+tmp[9464]*kernel[6]+tmp[9465]*kernel[7]+tmp[9466]*kernel[8];
				ans[9366]<=tmp[9265]*kernel[0]+tmp[9266]*kernel[1]+tmp[9267]*kernel[2]+tmp[9365]*kernel[3]+tmp[9366]*kernel[4]+tmp[9367]*kernel[5]+tmp[9465]*kernel[6]+tmp[9466]*kernel[7]+tmp[9467]*kernel[8];
				ans[9367]<=tmp[9266]*kernel[0]+tmp[9267]*kernel[1]+tmp[9268]*kernel[2]+tmp[9366]*kernel[3]+tmp[9367]*kernel[4]+tmp[9368]*kernel[5]+tmp[9466]*kernel[6]+tmp[9467]*kernel[7]+tmp[9468]*kernel[8];
				ans[9368]<=tmp[9267]*kernel[0]+tmp[9268]*kernel[1]+tmp[9269]*kernel[2]+tmp[9367]*kernel[3]+tmp[9368]*kernel[4]+tmp[9369]*kernel[5]+tmp[9467]*kernel[6]+tmp[9468]*kernel[7]+tmp[9469]*kernel[8];
				ans[9369]<=tmp[9268]*kernel[0]+tmp[9269]*kernel[1]+tmp[9270]*kernel[2]+tmp[9368]*kernel[3]+tmp[9369]*kernel[4]+tmp[9370]*kernel[5]+tmp[9468]*kernel[6]+tmp[9469]*kernel[7]+tmp[9470]*kernel[8];
				ans[9370]<=tmp[9269]*kernel[0]+tmp[9270]*kernel[1]+tmp[9271]*kernel[2]+tmp[9369]*kernel[3]+tmp[9370]*kernel[4]+tmp[9371]*kernel[5]+tmp[9469]*kernel[6]+tmp[9470]*kernel[7]+tmp[9471]*kernel[8];
				ans[9371]<=tmp[9270]*kernel[0]+tmp[9271]*kernel[1]+tmp[9272]*kernel[2]+tmp[9370]*kernel[3]+tmp[9371]*kernel[4]+tmp[9372]*kernel[5]+tmp[9470]*kernel[6]+tmp[9471]*kernel[7]+tmp[9472]*kernel[8];
				ans[9372]<=tmp[9271]*kernel[0]+tmp[9272]*kernel[1]+tmp[9273]*kernel[2]+tmp[9371]*kernel[3]+tmp[9372]*kernel[4]+tmp[9373]*kernel[5]+tmp[9471]*kernel[6]+tmp[9472]*kernel[7]+tmp[9473]*kernel[8];
				ans[9373]<=tmp[9272]*kernel[0]+tmp[9273]*kernel[1]+tmp[9274]*kernel[2]+tmp[9372]*kernel[3]+tmp[9373]*kernel[4]+tmp[9374]*kernel[5]+tmp[9472]*kernel[6]+tmp[9473]*kernel[7]+tmp[9474]*kernel[8];
				ans[9374]<=tmp[9273]*kernel[0]+tmp[9274]*kernel[1]+tmp[9275]*kernel[2]+tmp[9373]*kernel[3]+tmp[9374]*kernel[4]+tmp[9375]*kernel[5]+tmp[9473]*kernel[6]+tmp[9474]*kernel[7]+tmp[9475]*kernel[8];
				ans[9375]<=tmp[9274]*kernel[0]+tmp[9275]*kernel[1]+tmp[9276]*kernel[2]+tmp[9374]*kernel[3]+tmp[9375]*kernel[4]+tmp[9376]*kernel[5]+tmp[9474]*kernel[6]+tmp[9475]*kernel[7]+tmp[9476]*kernel[8];
				ans[9376]<=tmp[9275]*kernel[0]+tmp[9276]*kernel[1]+tmp[9277]*kernel[2]+tmp[9375]*kernel[3]+tmp[9376]*kernel[4]+tmp[9377]*kernel[5]+tmp[9475]*kernel[6]+tmp[9476]*kernel[7]+tmp[9477]*kernel[8];
				ans[9377]<=tmp[9276]*kernel[0]+tmp[9277]*kernel[1]+tmp[9278]*kernel[2]+tmp[9376]*kernel[3]+tmp[9377]*kernel[4]+tmp[9378]*kernel[5]+tmp[9476]*kernel[6]+tmp[9477]*kernel[7]+tmp[9478]*kernel[8];
				ans[9378]<=tmp[9277]*kernel[0]+tmp[9278]*kernel[1]+tmp[9279]*kernel[2]+tmp[9377]*kernel[3]+tmp[9378]*kernel[4]+tmp[9379]*kernel[5]+tmp[9477]*kernel[6]+tmp[9478]*kernel[7]+tmp[9479]*kernel[8];
				ans[9379]<=tmp[9278]*kernel[0]+tmp[9279]*kernel[1]+tmp[9280]*kernel[2]+tmp[9378]*kernel[3]+tmp[9379]*kernel[4]+tmp[9380]*kernel[5]+tmp[9478]*kernel[6]+tmp[9479]*kernel[7]+tmp[9480]*kernel[8];
				ans[9380]<=tmp[9279]*kernel[0]+tmp[9280]*kernel[1]+tmp[9281]*kernel[2]+tmp[9379]*kernel[3]+tmp[9380]*kernel[4]+tmp[9381]*kernel[5]+tmp[9479]*kernel[6]+tmp[9480]*kernel[7]+tmp[9481]*kernel[8];
				ans[9381]<=tmp[9280]*kernel[0]+tmp[9281]*kernel[1]+tmp[9282]*kernel[2]+tmp[9380]*kernel[3]+tmp[9381]*kernel[4]+tmp[9382]*kernel[5]+tmp[9480]*kernel[6]+tmp[9481]*kernel[7]+tmp[9482]*kernel[8];
				ans[9382]<=tmp[9281]*kernel[0]+tmp[9282]*kernel[1]+tmp[9283]*kernel[2]+tmp[9381]*kernel[3]+tmp[9382]*kernel[4]+tmp[9383]*kernel[5]+tmp[9481]*kernel[6]+tmp[9482]*kernel[7]+tmp[9483]*kernel[8];
				ans[9383]<=tmp[9282]*kernel[0]+tmp[9283]*kernel[1]+tmp[9284]*kernel[2]+tmp[9382]*kernel[3]+tmp[9383]*kernel[4]+tmp[9384]*kernel[5]+tmp[9482]*kernel[6]+tmp[9483]*kernel[7]+tmp[9484]*kernel[8];
				ans[9384]<=tmp[9283]*kernel[0]+tmp[9284]*kernel[1]+tmp[9285]*kernel[2]+tmp[9383]*kernel[3]+tmp[9384]*kernel[4]+tmp[9385]*kernel[5]+tmp[9483]*kernel[6]+tmp[9484]*kernel[7]+tmp[9485]*kernel[8];
				ans[9385]<=tmp[9284]*kernel[0]+tmp[9285]*kernel[1]+tmp[9286]*kernel[2]+tmp[9384]*kernel[3]+tmp[9385]*kernel[4]+tmp[9386]*kernel[5]+tmp[9484]*kernel[6]+tmp[9485]*kernel[7]+tmp[9486]*kernel[8];
				ans[9386]<=tmp[9285]*kernel[0]+tmp[9286]*kernel[1]+tmp[9287]*kernel[2]+tmp[9385]*kernel[3]+tmp[9386]*kernel[4]+tmp[9387]*kernel[5]+tmp[9485]*kernel[6]+tmp[9486]*kernel[7]+tmp[9487]*kernel[8];
				ans[9387]<=tmp[9286]*kernel[0]+tmp[9287]*kernel[1]+tmp[9288]*kernel[2]+tmp[9386]*kernel[3]+tmp[9387]*kernel[4]+tmp[9388]*kernel[5]+tmp[9486]*kernel[6]+tmp[9487]*kernel[7]+tmp[9488]*kernel[8];
				ans[9388]<=tmp[9287]*kernel[0]+tmp[9288]*kernel[1]+tmp[9289]*kernel[2]+tmp[9387]*kernel[3]+tmp[9388]*kernel[4]+tmp[9389]*kernel[5]+tmp[9487]*kernel[6]+tmp[9488]*kernel[7]+tmp[9489]*kernel[8];
				ans[9389]<=tmp[9288]*kernel[0]+tmp[9289]*kernel[1]+tmp[9290]*kernel[2]+tmp[9388]*kernel[3]+tmp[9389]*kernel[4]+tmp[9390]*kernel[5]+tmp[9488]*kernel[6]+tmp[9489]*kernel[7]+tmp[9490]*kernel[8];
				ans[9390]<=tmp[9289]*kernel[0]+tmp[9290]*kernel[1]+tmp[9291]*kernel[2]+tmp[9389]*kernel[3]+tmp[9390]*kernel[4]+tmp[9391]*kernel[5]+tmp[9489]*kernel[6]+tmp[9490]*kernel[7]+tmp[9491]*kernel[8];
				ans[9391]<=tmp[9290]*kernel[0]+tmp[9291]*kernel[1]+tmp[9292]*kernel[2]+tmp[9390]*kernel[3]+tmp[9391]*kernel[4]+tmp[9392]*kernel[5]+tmp[9490]*kernel[6]+tmp[9491]*kernel[7]+tmp[9492]*kernel[8];
				ans[9392]<=tmp[9291]*kernel[0]+tmp[9292]*kernel[1]+tmp[9293]*kernel[2]+tmp[9391]*kernel[3]+tmp[9392]*kernel[4]+tmp[9393]*kernel[5]+tmp[9491]*kernel[6]+tmp[9492]*kernel[7]+tmp[9493]*kernel[8];
				ans[9393]<=tmp[9292]*kernel[0]+tmp[9293]*kernel[1]+tmp[9294]*kernel[2]+tmp[9392]*kernel[3]+tmp[9393]*kernel[4]+tmp[9394]*kernel[5]+tmp[9492]*kernel[6]+tmp[9493]*kernel[7]+tmp[9494]*kernel[8];
				ans[9394]<=tmp[9293]*kernel[0]+tmp[9294]*kernel[1]+tmp[9295]*kernel[2]+tmp[9393]*kernel[3]+tmp[9394]*kernel[4]+tmp[9395]*kernel[5]+tmp[9493]*kernel[6]+tmp[9494]*kernel[7]+tmp[9495]*kernel[8];
				ans[9395]<=tmp[9294]*kernel[0]+tmp[9295]*kernel[1]+tmp[9296]*kernel[2]+tmp[9394]*kernel[3]+tmp[9395]*kernel[4]+tmp[9396]*kernel[5]+tmp[9494]*kernel[6]+tmp[9495]*kernel[7]+tmp[9496]*kernel[8];
				ans[9396]<=tmp[9295]*kernel[0]+tmp[9296]*kernel[1]+tmp[9297]*kernel[2]+tmp[9395]*kernel[3]+tmp[9396]*kernel[4]+tmp[9397]*kernel[5]+tmp[9495]*kernel[6]+tmp[9496]*kernel[7]+tmp[9497]*kernel[8];
				ans[9397]<=tmp[9296]*kernel[0]+tmp[9297]*kernel[1]+tmp[9298]*kernel[2]+tmp[9396]*kernel[3]+tmp[9397]*kernel[4]+tmp[9398]*kernel[5]+tmp[9496]*kernel[6]+tmp[9497]*kernel[7]+tmp[9498]*kernel[8];
				ans[9398]<=tmp[9297]*kernel[0]+tmp[9298]*kernel[1]+tmp[9299]*kernel[2]+tmp[9397]*kernel[3]+tmp[9398]*kernel[4]+tmp[9399]*kernel[5]+tmp[9497]*kernel[6]+tmp[9498]*kernel[7]+tmp[9499]*kernel[8];
				ans[9399]<=tmp[9298]*kernel[0]+tmp[9299]*kernel[1]+tmp[9398]*kernel[3]+tmp[9399]*kernel[4]+tmp[9498]*kernel[6]+tmp[9499]*kernel[7];
				ans[9400]<=tmp[9300]*kernel[1]+tmp[9301]*kernel[2]+tmp[9400]*kernel[4]+tmp[9401]*kernel[5]+tmp[9500]*kernel[7]+tmp[9501]*kernel[8];
				ans[9401]<=tmp[9300]*kernel[0]+tmp[9301]*kernel[1]+tmp[9302]*kernel[2]+tmp[9400]*kernel[3]+tmp[9401]*kernel[4]+tmp[9402]*kernel[5]+tmp[9500]*kernel[6]+tmp[9501]*kernel[7]+tmp[9502]*kernel[8];
				ans[9402]<=tmp[9301]*kernel[0]+tmp[9302]*kernel[1]+tmp[9303]*kernel[2]+tmp[9401]*kernel[3]+tmp[9402]*kernel[4]+tmp[9403]*kernel[5]+tmp[9501]*kernel[6]+tmp[9502]*kernel[7]+tmp[9503]*kernel[8];
				ans[9403]<=tmp[9302]*kernel[0]+tmp[9303]*kernel[1]+tmp[9304]*kernel[2]+tmp[9402]*kernel[3]+tmp[9403]*kernel[4]+tmp[9404]*kernel[5]+tmp[9502]*kernel[6]+tmp[9503]*kernel[7]+tmp[9504]*kernel[8];
				ans[9404]<=tmp[9303]*kernel[0]+tmp[9304]*kernel[1]+tmp[9305]*kernel[2]+tmp[9403]*kernel[3]+tmp[9404]*kernel[4]+tmp[9405]*kernel[5]+tmp[9503]*kernel[6]+tmp[9504]*kernel[7]+tmp[9505]*kernel[8];
				ans[9405]<=tmp[9304]*kernel[0]+tmp[9305]*kernel[1]+tmp[9306]*kernel[2]+tmp[9404]*kernel[3]+tmp[9405]*kernel[4]+tmp[9406]*kernel[5]+tmp[9504]*kernel[6]+tmp[9505]*kernel[7]+tmp[9506]*kernel[8];
				ans[9406]<=tmp[9305]*kernel[0]+tmp[9306]*kernel[1]+tmp[9307]*kernel[2]+tmp[9405]*kernel[3]+tmp[9406]*kernel[4]+tmp[9407]*kernel[5]+tmp[9505]*kernel[6]+tmp[9506]*kernel[7]+tmp[9507]*kernel[8];
				ans[9407]<=tmp[9306]*kernel[0]+tmp[9307]*kernel[1]+tmp[9308]*kernel[2]+tmp[9406]*kernel[3]+tmp[9407]*kernel[4]+tmp[9408]*kernel[5]+tmp[9506]*kernel[6]+tmp[9507]*kernel[7]+tmp[9508]*kernel[8];
				ans[9408]<=tmp[9307]*kernel[0]+tmp[9308]*kernel[1]+tmp[9309]*kernel[2]+tmp[9407]*kernel[3]+tmp[9408]*kernel[4]+tmp[9409]*kernel[5]+tmp[9507]*kernel[6]+tmp[9508]*kernel[7]+tmp[9509]*kernel[8];
				ans[9409]<=tmp[9308]*kernel[0]+tmp[9309]*kernel[1]+tmp[9310]*kernel[2]+tmp[9408]*kernel[3]+tmp[9409]*kernel[4]+tmp[9410]*kernel[5]+tmp[9508]*kernel[6]+tmp[9509]*kernel[7]+tmp[9510]*kernel[8];
				ans[9410]<=tmp[9309]*kernel[0]+tmp[9310]*kernel[1]+tmp[9311]*kernel[2]+tmp[9409]*kernel[3]+tmp[9410]*kernel[4]+tmp[9411]*kernel[5]+tmp[9509]*kernel[6]+tmp[9510]*kernel[7]+tmp[9511]*kernel[8];
				ans[9411]<=tmp[9310]*kernel[0]+tmp[9311]*kernel[1]+tmp[9312]*kernel[2]+tmp[9410]*kernel[3]+tmp[9411]*kernel[4]+tmp[9412]*kernel[5]+tmp[9510]*kernel[6]+tmp[9511]*kernel[7]+tmp[9512]*kernel[8];
				ans[9412]<=tmp[9311]*kernel[0]+tmp[9312]*kernel[1]+tmp[9313]*kernel[2]+tmp[9411]*kernel[3]+tmp[9412]*kernel[4]+tmp[9413]*kernel[5]+tmp[9511]*kernel[6]+tmp[9512]*kernel[7]+tmp[9513]*kernel[8];
				ans[9413]<=tmp[9312]*kernel[0]+tmp[9313]*kernel[1]+tmp[9314]*kernel[2]+tmp[9412]*kernel[3]+tmp[9413]*kernel[4]+tmp[9414]*kernel[5]+tmp[9512]*kernel[6]+tmp[9513]*kernel[7]+tmp[9514]*kernel[8];
				ans[9414]<=tmp[9313]*kernel[0]+tmp[9314]*kernel[1]+tmp[9315]*kernel[2]+tmp[9413]*kernel[3]+tmp[9414]*kernel[4]+tmp[9415]*kernel[5]+tmp[9513]*kernel[6]+tmp[9514]*kernel[7]+tmp[9515]*kernel[8];
				ans[9415]<=tmp[9314]*kernel[0]+tmp[9315]*kernel[1]+tmp[9316]*kernel[2]+tmp[9414]*kernel[3]+tmp[9415]*kernel[4]+tmp[9416]*kernel[5]+tmp[9514]*kernel[6]+tmp[9515]*kernel[7]+tmp[9516]*kernel[8];
				ans[9416]<=tmp[9315]*kernel[0]+tmp[9316]*kernel[1]+tmp[9317]*kernel[2]+tmp[9415]*kernel[3]+tmp[9416]*kernel[4]+tmp[9417]*kernel[5]+tmp[9515]*kernel[6]+tmp[9516]*kernel[7]+tmp[9517]*kernel[8];
				ans[9417]<=tmp[9316]*kernel[0]+tmp[9317]*kernel[1]+tmp[9318]*kernel[2]+tmp[9416]*kernel[3]+tmp[9417]*kernel[4]+tmp[9418]*kernel[5]+tmp[9516]*kernel[6]+tmp[9517]*kernel[7]+tmp[9518]*kernel[8];
				ans[9418]<=tmp[9317]*kernel[0]+tmp[9318]*kernel[1]+tmp[9319]*kernel[2]+tmp[9417]*kernel[3]+tmp[9418]*kernel[4]+tmp[9419]*kernel[5]+tmp[9517]*kernel[6]+tmp[9518]*kernel[7]+tmp[9519]*kernel[8];
				ans[9419]<=tmp[9318]*kernel[0]+tmp[9319]*kernel[1]+tmp[9320]*kernel[2]+tmp[9418]*kernel[3]+tmp[9419]*kernel[4]+tmp[9420]*kernel[5]+tmp[9518]*kernel[6]+tmp[9519]*kernel[7]+tmp[9520]*kernel[8];
				ans[9420]<=tmp[9319]*kernel[0]+tmp[9320]*kernel[1]+tmp[9321]*kernel[2]+tmp[9419]*kernel[3]+tmp[9420]*kernel[4]+tmp[9421]*kernel[5]+tmp[9519]*kernel[6]+tmp[9520]*kernel[7]+tmp[9521]*kernel[8];
				ans[9421]<=tmp[9320]*kernel[0]+tmp[9321]*kernel[1]+tmp[9322]*kernel[2]+tmp[9420]*kernel[3]+tmp[9421]*kernel[4]+tmp[9422]*kernel[5]+tmp[9520]*kernel[6]+tmp[9521]*kernel[7]+tmp[9522]*kernel[8];
				ans[9422]<=tmp[9321]*kernel[0]+tmp[9322]*kernel[1]+tmp[9323]*kernel[2]+tmp[9421]*kernel[3]+tmp[9422]*kernel[4]+tmp[9423]*kernel[5]+tmp[9521]*kernel[6]+tmp[9522]*kernel[7]+tmp[9523]*kernel[8];
				ans[9423]<=tmp[9322]*kernel[0]+tmp[9323]*kernel[1]+tmp[9324]*kernel[2]+tmp[9422]*kernel[3]+tmp[9423]*kernel[4]+tmp[9424]*kernel[5]+tmp[9522]*kernel[6]+tmp[9523]*kernel[7]+tmp[9524]*kernel[8];
				ans[9424]<=tmp[9323]*kernel[0]+tmp[9324]*kernel[1]+tmp[9325]*kernel[2]+tmp[9423]*kernel[3]+tmp[9424]*kernel[4]+tmp[9425]*kernel[5]+tmp[9523]*kernel[6]+tmp[9524]*kernel[7]+tmp[9525]*kernel[8];
				ans[9425]<=tmp[9324]*kernel[0]+tmp[9325]*kernel[1]+tmp[9326]*kernel[2]+tmp[9424]*kernel[3]+tmp[9425]*kernel[4]+tmp[9426]*kernel[5]+tmp[9524]*kernel[6]+tmp[9525]*kernel[7]+tmp[9526]*kernel[8];
				ans[9426]<=tmp[9325]*kernel[0]+tmp[9326]*kernel[1]+tmp[9327]*kernel[2]+tmp[9425]*kernel[3]+tmp[9426]*kernel[4]+tmp[9427]*kernel[5]+tmp[9525]*kernel[6]+tmp[9526]*kernel[7]+tmp[9527]*kernel[8];
				ans[9427]<=tmp[9326]*kernel[0]+tmp[9327]*kernel[1]+tmp[9328]*kernel[2]+tmp[9426]*kernel[3]+tmp[9427]*kernel[4]+tmp[9428]*kernel[5]+tmp[9526]*kernel[6]+tmp[9527]*kernel[7]+tmp[9528]*kernel[8];
				ans[9428]<=tmp[9327]*kernel[0]+tmp[9328]*kernel[1]+tmp[9329]*kernel[2]+tmp[9427]*kernel[3]+tmp[9428]*kernel[4]+tmp[9429]*kernel[5]+tmp[9527]*kernel[6]+tmp[9528]*kernel[7]+tmp[9529]*kernel[8];
				ans[9429]<=tmp[9328]*kernel[0]+tmp[9329]*kernel[1]+tmp[9330]*kernel[2]+tmp[9428]*kernel[3]+tmp[9429]*kernel[4]+tmp[9430]*kernel[5]+tmp[9528]*kernel[6]+tmp[9529]*kernel[7]+tmp[9530]*kernel[8];
				ans[9430]<=tmp[9329]*kernel[0]+tmp[9330]*kernel[1]+tmp[9331]*kernel[2]+tmp[9429]*kernel[3]+tmp[9430]*kernel[4]+tmp[9431]*kernel[5]+tmp[9529]*kernel[6]+tmp[9530]*kernel[7]+tmp[9531]*kernel[8];
				ans[9431]<=tmp[9330]*kernel[0]+tmp[9331]*kernel[1]+tmp[9332]*kernel[2]+tmp[9430]*kernel[3]+tmp[9431]*kernel[4]+tmp[9432]*kernel[5]+tmp[9530]*kernel[6]+tmp[9531]*kernel[7]+tmp[9532]*kernel[8];
				ans[9432]<=tmp[9331]*kernel[0]+tmp[9332]*kernel[1]+tmp[9333]*kernel[2]+tmp[9431]*kernel[3]+tmp[9432]*kernel[4]+tmp[9433]*kernel[5]+tmp[9531]*kernel[6]+tmp[9532]*kernel[7]+tmp[9533]*kernel[8];
				ans[9433]<=tmp[9332]*kernel[0]+tmp[9333]*kernel[1]+tmp[9334]*kernel[2]+tmp[9432]*kernel[3]+tmp[9433]*kernel[4]+tmp[9434]*kernel[5]+tmp[9532]*kernel[6]+tmp[9533]*kernel[7]+tmp[9534]*kernel[8];
				ans[9434]<=tmp[9333]*kernel[0]+tmp[9334]*kernel[1]+tmp[9335]*kernel[2]+tmp[9433]*kernel[3]+tmp[9434]*kernel[4]+tmp[9435]*kernel[5]+tmp[9533]*kernel[6]+tmp[9534]*kernel[7]+tmp[9535]*kernel[8];
				ans[9435]<=tmp[9334]*kernel[0]+tmp[9335]*kernel[1]+tmp[9336]*kernel[2]+tmp[9434]*kernel[3]+tmp[9435]*kernel[4]+tmp[9436]*kernel[5]+tmp[9534]*kernel[6]+tmp[9535]*kernel[7]+tmp[9536]*kernel[8];
				ans[9436]<=tmp[9335]*kernel[0]+tmp[9336]*kernel[1]+tmp[9337]*kernel[2]+tmp[9435]*kernel[3]+tmp[9436]*kernel[4]+tmp[9437]*kernel[5]+tmp[9535]*kernel[6]+tmp[9536]*kernel[7]+tmp[9537]*kernel[8];
				ans[9437]<=tmp[9336]*kernel[0]+tmp[9337]*kernel[1]+tmp[9338]*kernel[2]+tmp[9436]*kernel[3]+tmp[9437]*kernel[4]+tmp[9438]*kernel[5]+tmp[9536]*kernel[6]+tmp[9537]*kernel[7]+tmp[9538]*kernel[8];
				ans[9438]<=tmp[9337]*kernel[0]+tmp[9338]*kernel[1]+tmp[9339]*kernel[2]+tmp[9437]*kernel[3]+tmp[9438]*kernel[4]+tmp[9439]*kernel[5]+tmp[9537]*kernel[6]+tmp[9538]*kernel[7]+tmp[9539]*kernel[8];
				ans[9439]<=tmp[9338]*kernel[0]+tmp[9339]*kernel[1]+tmp[9340]*kernel[2]+tmp[9438]*kernel[3]+tmp[9439]*kernel[4]+tmp[9440]*kernel[5]+tmp[9538]*kernel[6]+tmp[9539]*kernel[7]+tmp[9540]*kernel[8];
				ans[9440]<=tmp[9339]*kernel[0]+tmp[9340]*kernel[1]+tmp[9341]*kernel[2]+tmp[9439]*kernel[3]+tmp[9440]*kernel[4]+tmp[9441]*kernel[5]+tmp[9539]*kernel[6]+tmp[9540]*kernel[7]+tmp[9541]*kernel[8];
				ans[9441]<=tmp[9340]*kernel[0]+tmp[9341]*kernel[1]+tmp[9342]*kernel[2]+tmp[9440]*kernel[3]+tmp[9441]*kernel[4]+tmp[9442]*kernel[5]+tmp[9540]*kernel[6]+tmp[9541]*kernel[7]+tmp[9542]*kernel[8];
				ans[9442]<=tmp[9341]*kernel[0]+tmp[9342]*kernel[1]+tmp[9343]*kernel[2]+tmp[9441]*kernel[3]+tmp[9442]*kernel[4]+tmp[9443]*kernel[5]+tmp[9541]*kernel[6]+tmp[9542]*kernel[7]+tmp[9543]*kernel[8];
				ans[9443]<=tmp[9342]*kernel[0]+tmp[9343]*kernel[1]+tmp[9344]*kernel[2]+tmp[9442]*kernel[3]+tmp[9443]*kernel[4]+tmp[9444]*kernel[5]+tmp[9542]*kernel[6]+tmp[9543]*kernel[7]+tmp[9544]*kernel[8];
				ans[9444]<=tmp[9343]*kernel[0]+tmp[9344]*kernel[1]+tmp[9345]*kernel[2]+tmp[9443]*kernel[3]+tmp[9444]*kernel[4]+tmp[9445]*kernel[5]+tmp[9543]*kernel[6]+tmp[9544]*kernel[7]+tmp[9545]*kernel[8];
				ans[9445]<=tmp[9344]*kernel[0]+tmp[9345]*kernel[1]+tmp[9346]*kernel[2]+tmp[9444]*kernel[3]+tmp[9445]*kernel[4]+tmp[9446]*kernel[5]+tmp[9544]*kernel[6]+tmp[9545]*kernel[7]+tmp[9546]*kernel[8];
				ans[9446]<=tmp[9345]*kernel[0]+tmp[9346]*kernel[1]+tmp[9347]*kernel[2]+tmp[9445]*kernel[3]+tmp[9446]*kernel[4]+tmp[9447]*kernel[5]+tmp[9545]*kernel[6]+tmp[9546]*kernel[7]+tmp[9547]*kernel[8];
				ans[9447]<=tmp[9346]*kernel[0]+tmp[9347]*kernel[1]+tmp[9348]*kernel[2]+tmp[9446]*kernel[3]+tmp[9447]*kernel[4]+tmp[9448]*kernel[5]+tmp[9546]*kernel[6]+tmp[9547]*kernel[7]+tmp[9548]*kernel[8];
				ans[9448]<=tmp[9347]*kernel[0]+tmp[9348]*kernel[1]+tmp[9349]*kernel[2]+tmp[9447]*kernel[3]+tmp[9448]*kernel[4]+tmp[9449]*kernel[5]+tmp[9547]*kernel[6]+tmp[9548]*kernel[7]+tmp[9549]*kernel[8];
				ans[9449]<=tmp[9348]*kernel[0]+tmp[9349]*kernel[1]+tmp[9350]*kernel[2]+tmp[9448]*kernel[3]+tmp[9449]*kernel[4]+tmp[9450]*kernel[5]+tmp[9548]*kernel[6]+tmp[9549]*kernel[7]+tmp[9550]*kernel[8];
				ans[9450]<=tmp[9349]*kernel[0]+tmp[9350]*kernel[1]+tmp[9351]*kernel[2]+tmp[9449]*kernel[3]+tmp[9450]*kernel[4]+tmp[9451]*kernel[5]+tmp[9549]*kernel[6]+tmp[9550]*kernel[7]+tmp[9551]*kernel[8];
				ans[9451]<=tmp[9350]*kernel[0]+tmp[9351]*kernel[1]+tmp[9352]*kernel[2]+tmp[9450]*kernel[3]+tmp[9451]*kernel[4]+tmp[9452]*kernel[5]+tmp[9550]*kernel[6]+tmp[9551]*kernel[7]+tmp[9552]*kernel[8];
				ans[9452]<=tmp[9351]*kernel[0]+tmp[9352]*kernel[1]+tmp[9353]*kernel[2]+tmp[9451]*kernel[3]+tmp[9452]*kernel[4]+tmp[9453]*kernel[5]+tmp[9551]*kernel[6]+tmp[9552]*kernel[7]+tmp[9553]*kernel[8];
				ans[9453]<=tmp[9352]*kernel[0]+tmp[9353]*kernel[1]+tmp[9354]*kernel[2]+tmp[9452]*kernel[3]+tmp[9453]*kernel[4]+tmp[9454]*kernel[5]+tmp[9552]*kernel[6]+tmp[9553]*kernel[7]+tmp[9554]*kernel[8];
				ans[9454]<=tmp[9353]*kernel[0]+tmp[9354]*kernel[1]+tmp[9355]*kernel[2]+tmp[9453]*kernel[3]+tmp[9454]*kernel[4]+tmp[9455]*kernel[5]+tmp[9553]*kernel[6]+tmp[9554]*kernel[7]+tmp[9555]*kernel[8];
				ans[9455]<=tmp[9354]*kernel[0]+tmp[9355]*kernel[1]+tmp[9356]*kernel[2]+tmp[9454]*kernel[3]+tmp[9455]*kernel[4]+tmp[9456]*kernel[5]+tmp[9554]*kernel[6]+tmp[9555]*kernel[7]+tmp[9556]*kernel[8];
				ans[9456]<=tmp[9355]*kernel[0]+tmp[9356]*kernel[1]+tmp[9357]*kernel[2]+tmp[9455]*kernel[3]+tmp[9456]*kernel[4]+tmp[9457]*kernel[5]+tmp[9555]*kernel[6]+tmp[9556]*kernel[7]+tmp[9557]*kernel[8];
				ans[9457]<=tmp[9356]*kernel[0]+tmp[9357]*kernel[1]+tmp[9358]*kernel[2]+tmp[9456]*kernel[3]+tmp[9457]*kernel[4]+tmp[9458]*kernel[5]+tmp[9556]*kernel[6]+tmp[9557]*kernel[7]+tmp[9558]*kernel[8];
				ans[9458]<=tmp[9357]*kernel[0]+tmp[9358]*kernel[1]+tmp[9359]*kernel[2]+tmp[9457]*kernel[3]+tmp[9458]*kernel[4]+tmp[9459]*kernel[5]+tmp[9557]*kernel[6]+tmp[9558]*kernel[7]+tmp[9559]*kernel[8];
				ans[9459]<=tmp[9358]*kernel[0]+tmp[9359]*kernel[1]+tmp[9360]*kernel[2]+tmp[9458]*kernel[3]+tmp[9459]*kernel[4]+tmp[9460]*kernel[5]+tmp[9558]*kernel[6]+tmp[9559]*kernel[7]+tmp[9560]*kernel[8];
				ans[9460]<=tmp[9359]*kernel[0]+tmp[9360]*kernel[1]+tmp[9361]*kernel[2]+tmp[9459]*kernel[3]+tmp[9460]*kernel[4]+tmp[9461]*kernel[5]+tmp[9559]*kernel[6]+tmp[9560]*kernel[7]+tmp[9561]*kernel[8];
				ans[9461]<=tmp[9360]*kernel[0]+tmp[9361]*kernel[1]+tmp[9362]*kernel[2]+tmp[9460]*kernel[3]+tmp[9461]*kernel[4]+tmp[9462]*kernel[5]+tmp[9560]*kernel[6]+tmp[9561]*kernel[7]+tmp[9562]*kernel[8];
				ans[9462]<=tmp[9361]*kernel[0]+tmp[9362]*kernel[1]+tmp[9363]*kernel[2]+tmp[9461]*kernel[3]+tmp[9462]*kernel[4]+tmp[9463]*kernel[5]+tmp[9561]*kernel[6]+tmp[9562]*kernel[7]+tmp[9563]*kernel[8];
				ans[9463]<=tmp[9362]*kernel[0]+tmp[9363]*kernel[1]+tmp[9364]*kernel[2]+tmp[9462]*kernel[3]+tmp[9463]*kernel[4]+tmp[9464]*kernel[5]+tmp[9562]*kernel[6]+tmp[9563]*kernel[7]+tmp[9564]*kernel[8];
				ans[9464]<=tmp[9363]*kernel[0]+tmp[9364]*kernel[1]+tmp[9365]*kernel[2]+tmp[9463]*kernel[3]+tmp[9464]*kernel[4]+tmp[9465]*kernel[5]+tmp[9563]*kernel[6]+tmp[9564]*kernel[7]+tmp[9565]*kernel[8];
				ans[9465]<=tmp[9364]*kernel[0]+tmp[9365]*kernel[1]+tmp[9366]*kernel[2]+tmp[9464]*kernel[3]+tmp[9465]*kernel[4]+tmp[9466]*kernel[5]+tmp[9564]*kernel[6]+tmp[9565]*kernel[7]+tmp[9566]*kernel[8];
				ans[9466]<=tmp[9365]*kernel[0]+tmp[9366]*kernel[1]+tmp[9367]*kernel[2]+tmp[9465]*kernel[3]+tmp[9466]*kernel[4]+tmp[9467]*kernel[5]+tmp[9565]*kernel[6]+tmp[9566]*kernel[7]+tmp[9567]*kernel[8];
				ans[9467]<=tmp[9366]*kernel[0]+tmp[9367]*kernel[1]+tmp[9368]*kernel[2]+tmp[9466]*kernel[3]+tmp[9467]*kernel[4]+tmp[9468]*kernel[5]+tmp[9566]*kernel[6]+tmp[9567]*kernel[7]+tmp[9568]*kernel[8];
				ans[9468]<=tmp[9367]*kernel[0]+tmp[9368]*kernel[1]+tmp[9369]*kernel[2]+tmp[9467]*kernel[3]+tmp[9468]*kernel[4]+tmp[9469]*kernel[5]+tmp[9567]*kernel[6]+tmp[9568]*kernel[7]+tmp[9569]*kernel[8];
				ans[9469]<=tmp[9368]*kernel[0]+tmp[9369]*kernel[1]+tmp[9370]*kernel[2]+tmp[9468]*kernel[3]+tmp[9469]*kernel[4]+tmp[9470]*kernel[5]+tmp[9568]*kernel[6]+tmp[9569]*kernel[7]+tmp[9570]*kernel[8];
				ans[9470]<=tmp[9369]*kernel[0]+tmp[9370]*kernel[1]+tmp[9371]*kernel[2]+tmp[9469]*kernel[3]+tmp[9470]*kernel[4]+tmp[9471]*kernel[5]+tmp[9569]*kernel[6]+tmp[9570]*kernel[7]+tmp[9571]*kernel[8];
				ans[9471]<=tmp[9370]*kernel[0]+tmp[9371]*kernel[1]+tmp[9372]*kernel[2]+tmp[9470]*kernel[3]+tmp[9471]*kernel[4]+tmp[9472]*kernel[5]+tmp[9570]*kernel[6]+tmp[9571]*kernel[7]+tmp[9572]*kernel[8];
				ans[9472]<=tmp[9371]*kernel[0]+tmp[9372]*kernel[1]+tmp[9373]*kernel[2]+tmp[9471]*kernel[3]+tmp[9472]*kernel[4]+tmp[9473]*kernel[5]+tmp[9571]*kernel[6]+tmp[9572]*kernel[7]+tmp[9573]*kernel[8];
				ans[9473]<=tmp[9372]*kernel[0]+tmp[9373]*kernel[1]+tmp[9374]*kernel[2]+tmp[9472]*kernel[3]+tmp[9473]*kernel[4]+tmp[9474]*kernel[5]+tmp[9572]*kernel[6]+tmp[9573]*kernel[7]+tmp[9574]*kernel[8];
				ans[9474]<=tmp[9373]*kernel[0]+tmp[9374]*kernel[1]+tmp[9375]*kernel[2]+tmp[9473]*kernel[3]+tmp[9474]*kernel[4]+tmp[9475]*kernel[5]+tmp[9573]*kernel[6]+tmp[9574]*kernel[7]+tmp[9575]*kernel[8];
				ans[9475]<=tmp[9374]*kernel[0]+tmp[9375]*kernel[1]+tmp[9376]*kernel[2]+tmp[9474]*kernel[3]+tmp[9475]*kernel[4]+tmp[9476]*kernel[5]+tmp[9574]*kernel[6]+tmp[9575]*kernel[7]+tmp[9576]*kernel[8];
				ans[9476]<=tmp[9375]*kernel[0]+tmp[9376]*kernel[1]+tmp[9377]*kernel[2]+tmp[9475]*kernel[3]+tmp[9476]*kernel[4]+tmp[9477]*kernel[5]+tmp[9575]*kernel[6]+tmp[9576]*kernel[7]+tmp[9577]*kernel[8];
				ans[9477]<=tmp[9376]*kernel[0]+tmp[9377]*kernel[1]+tmp[9378]*kernel[2]+tmp[9476]*kernel[3]+tmp[9477]*kernel[4]+tmp[9478]*kernel[5]+tmp[9576]*kernel[6]+tmp[9577]*kernel[7]+tmp[9578]*kernel[8];
				ans[9478]<=tmp[9377]*kernel[0]+tmp[9378]*kernel[1]+tmp[9379]*kernel[2]+tmp[9477]*kernel[3]+tmp[9478]*kernel[4]+tmp[9479]*kernel[5]+tmp[9577]*kernel[6]+tmp[9578]*kernel[7]+tmp[9579]*kernel[8];
				ans[9479]<=tmp[9378]*kernel[0]+tmp[9379]*kernel[1]+tmp[9380]*kernel[2]+tmp[9478]*kernel[3]+tmp[9479]*kernel[4]+tmp[9480]*kernel[5]+tmp[9578]*kernel[6]+tmp[9579]*kernel[7]+tmp[9580]*kernel[8];
				ans[9480]<=tmp[9379]*kernel[0]+tmp[9380]*kernel[1]+tmp[9381]*kernel[2]+tmp[9479]*kernel[3]+tmp[9480]*kernel[4]+tmp[9481]*kernel[5]+tmp[9579]*kernel[6]+tmp[9580]*kernel[7]+tmp[9581]*kernel[8];
				ans[9481]<=tmp[9380]*kernel[0]+tmp[9381]*kernel[1]+tmp[9382]*kernel[2]+tmp[9480]*kernel[3]+tmp[9481]*kernel[4]+tmp[9482]*kernel[5]+tmp[9580]*kernel[6]+tmp[9581]*kernel[7]+tmp[9582]*kernel[8];
				ans[9482]<=tmp[9381]*kernel[0]+tmp[9382]*kernel[1]+tmp[9383]*kernel[2]+tmp[9481]*kernel[3]+tmp[9482]*kernel[4]+tmp[9483]*kernel[5]+tmp[9581]*kernel[6]+tmp[9582]*kernel[7]+tmp[9583]*kernel[8];
				ans[9483]<=tmp[9382]*kernel[0]+tmp[9383]*kernel[1]+tmp[9384]*kernel[2]+tmp[9482]*kernel[3]+tmp[9483]*kernel[4]+tmp[9484]*kernel[5]+tmp[9582]*kernel[6]+tmp[9583]*kernel[7]+tmp[9584]*kernel[8];
				ans[9484]<=tmp[9383]*kernel[0]+tmp[9384]*kernel[1]+tmp[9385]*kernel[2]+tmp[9483]*kernel[3]+tmp[9484]*kernel[4]+tmp[9485]*kernel[5]+tmp[9583]*kernel[6]+tmp[9584]*kernel[7]+tmp[9585]*kernel[8];
				ans[9485]<=tmp[9384]*kernel[0]+tmp[9385]*kernel[1]+tmp[9386]*kernel[2]+tmp[9484]*kernel[3]+tmp[9485]*kernel[4]+tmp[9486]*kernel[5]+tmp[9584]*kernel[6]+tmp[9585]*kernel[7]+tmp[9586]*kernel[8];
				ans[9486]<=tmp[9385]*kernel[0]+tmp[9386]*kernel[1]+tmp[9387]*kernel[2]+tmp[9485]*kernel[3]+tmp[9486]*kernel[4]+tmp[9487]*kernel[5]+tmp[9585]*kernel[6]+tmp[9586]*kernel[7]+tmp[9587]*kernel[8];
				ans[9487]<=tmp[9386]*kernel[0]+tmp[9387]*kernel[1]+tmp[9388]*kernel[2]+tmp[9486]*kernel[3]+tmp[9487]*kernel[4]+tmp[9488]*kernel[5]+tmp[9586]*kernel[6]+tmp[9587]*kernel[7]+tmp[9588]*kernel[8];
				ans[9488]<=tmp[9387]*kernel[0]+tmp[9388]*kernel[1]+tmp[9389]*kernel[2]+tmp[9487]*kernel[3]+tmp[9488]*kernel[4]+tmp[9489]*kernel[5]+tmp[9587]*kernel[6]+tmp[9588]*kernel[7]+tmp[9589]*kernel[8];
				ans[9489]<=tmp[9388]*kernel[0]+tmp[9389]*kernel[1]+tmp[9390]*kernel[2]+tmp[9488]*kernel[3]+tmp[9489]*kernel[4]+tmp[9490]*kernel[5]+tmp[9588]*kernel[6]+tmp[9589]*kernel[7]+tmp[9590]*kernel[8];
				ans[9490]<=tmp[9389]*kernel[0]+tmp[9390]*kernel[1]+tmp[9391]*kernel[2]+tmp[9489]*kernel[3]+tmp[9490]*kernel[4]+tmp[9491]*kernel[5]+tmp[9589]*kernel[6]+tmp[9590]*kernel[7]+tmp[9591]*kernel[8];
				ans[9491]<=tmp[9390]*kernel[0]+tmp[9391]*kernel[1]+tmp[9392]*kernel[2]+tmp[9490]*kernel[3]+tmp[9491]*kernel[4]+tmp[9492]*kernel[5]+tmp[9590]*kernel[6]+tmp[9591]*kernel[7]+tmp[9592]*kernel[8];
				ans[9492]<=tmp[9391]*kernel[0]+tmp[9392]*kernel[1]+tmp[9393]*kernel[2]+tmp[9491]*kernel[3]+tmp[9492]*kernel[4]+tmp[9493]*kernel[5]+tmp[9591]*kernel[6]+tmp[9592]*kernel[7]+tmp[9593]*kernel[8];
				ans[9493]<=tmp[9392]*kernel[0]+tmp[9393]*kernel[1]+tmp[9394]*kernel[2]+tmp[9492]*kernel[3]+tmp[9493]*kernel[4]+tmp[9494]*kernel[5]+tmp[9592]*kernel[6]+tmp[9593]*kernel[7]+tmp[9594]*kernel[8];
				ans[9494]<=tmp[9393]*kernel[0]+tmp[9394]*kernel[1]+tmp[9395]*kernel[2]+tmp[9493]*kernel[3]+tmp[9494]*kernel[4]+tmp[9495]*kernel[5]+tmp[9593]*kernel[6]+tmp[9594]*kernel[7]+tmp[9595]*kernel[8];
				ans[9495]<=tmp[9394]*kernel[0]+tmp[9395]*kernel[1]+tmp[9396]*kernel[2]+tmp[9494]*kernel[3]+tmp[9495]*kernel[4]+tmp[9496]*kernel[5]+tmp[9594]*kernel[6]+tmp[9595]*kernel[7]+tmp[9596]*kernel[8];
				ans[9496]<=tmp[9395]*kernel[0]+tmp[9396]*kernel[1]+tmp[9397]*kernel[2]+tmp[9495]*kernel[3]+tmp[9496]*kernel[4]+tmp[9497]*kernel[5]+tmp[9595]*kernel[6]+tmp[9596]*kernel[7]+tmp[9597]*kernel[8];
				ans[9497]<=tmp[9396]*kernel[0]+tmp[9397]*kernel[1]+tmp[9398]*kernel[2]+tmp[9496]*kernel[3]+tmp[9497]*kernel[4]+tmp[9498]*kernel[5]+tmp[9596]*kernel[6]+tmp[9597]*kernel[7]+tmp[9598]*kernel[8];
				ans[9498]<=tmp[9397]*kernel[0]+tmp[9398]*kernel[1]+tmp[9399]*kernel[2]+tmp[9497]*kernel[3]+tmp[9498]*kernel[4]+tmp[9499]*kernel[5]+tmp[9597]*kernel[6]+tmp[9598]*kernel[7]+tmp[9599]*kernel[8];
				ans[9499]<=tmp[9398]*kernel[0]+tmp[9399]*kernel[1]+tmp[9498]*kernel[3]+tmp[9499]*kernel[4]+tmp[9598]*kernel[6]+tmp[9599]*kernel[7];
				ans[9500]<=tmp[9400]*kernel[1]+tmp[9401]*kernel[2]+tmp[9500]*kernel[4]+tmp[9501]*kernel[5]+tmp[9600]*kernel[7]+tmp[9601]*kernel[8];
				ans[9501]<=tmp[9400]*kernel[0]+tmp[9401]*kernel[1]+tmp[9402]*kernel[2]+tmp[9500]*kernel[3]+tmp[9501]*kernel[4]+tmp[9502]*kernel[5]+tmp[9600]*kernel[6]+tmp[9601]*kernel[7]+tmp[9602]*kernel[8];
				ans[9502]<=tmp[9401]*kernel[0]+tmp[9402]*kernel[1]+tmp[9403]*kernel[2]+tmp[9501]*kernel[3]+tmp[9502]*kernel[4]+tmp[9503]*kernel[5]+tmp[9601]*kernel[6]+tmp[9602]*kernel[7]+tmp[9603]*kernel[8];
				ans[9503]<=tmp[9402]*kernel[0]+tmp[9403]*kernel[1]+tmp[9404]*kernel[2]+tmp[9502]*kernel[3]+tmp[9503]*kernel[4]+tmp[9504]*kernel[5]+tmp[9602]*kernel[6]+tmp[9603]*kernel[7]+tmp[9604]*kernel[8];
				ans[9504]<=tmp[9403]*kernel[0]+tmp[9404]*kernel[1]+tmp[9405]*kernel[2]+tmp[9503]*kernel[3]+tmp[9504]*kernel[4]+tmp[9505]*kernel[5]+tmp[9603]*kernel[6]+tmp[9604]*kernel[7]+tmp[9605]*kernel[8];
				ans[9505]<=tmp[9404]*kernel[0]+tmp[9405]*kernel[1]+tmp[9406]*kernel[2]+tmp[9504]*kernel[3]+tmp[9505]*kernel[4]+tmp[9506]*kernel[5]+tmp[9604]*kernel[6]+tmp[9605]*kernel[7]+tmp[9606]*kernel[8];
				ans[9506]<=tmp[9405]*kernel[0]+tmp[9406]*kernel[1]+tmp[9407]*kernel[2]+tmp[9505]*kernel[3]+tmp[9506]*kernel[4]+tmp[9507]*kernel[5]+tmp[9605]*kernel[6]+tmp[9606]*kernel[7]+tmp[9607]*kernel[8];
				ans[9507]<=tmp[9406]*kernel[0]+tmp[9407]*kernel[1]+tmp[9408]*kernel[2]+tmp[9506]*kernel[3]+tmp[9507]*kernel[4]+tmp[9508]*kernel[5]+tmp[9606]*kernel[6]+tmp[9607]*kernel[7]+tmp[9608]*kernel[8];
				ans[9508]<=tmp[9407]*kernel[0]+tmp[9408]*kernel[1]+tmp[9409]*kernel[2]+tmp[9507]*kernel[3]+tmp[9508]*kernel[4]+tmp[9509]*kernel[5]+tmp[9607]*kernel[6]+tmp[9608]*kernel[7]+tmp[9609]*kernel[8];
				ans[9509]<=tmp[9408]*kernel[0]+tmp[9409]*kernel[1]+tmp[9410]*kernel[2]+tmp[9508]*kernel[3]+tmp[9509]*kernel[4]+tmp[9510]*kernel[5]+tmp[9608]*kernel[6]+tmp[9609]*kernel[7]+tmp[9610]*kernel[8];
				ans[9510]<=tmp[9409]*kernel[0]+tmp[9410]*kernel[1]+tmp[9411]*kernel[2]+tmp[9509]*kernel[3]+tmp[9510]*kernel[4]+tmp[9511]*kernel[5]+tmp[9609]*kernel[6]+tmp[9610]*kernel[7]+tmp[9611]*kernel[8];
				ans[9511]<=tmp[9410]*kernel[0]+tmp[9411]*kernel[1]+tmp[9412]*kernel[2]+tmp[9510]*kernel[3]+tmp[9511]*kernel[4]+tmp[9512]*kernel[5]+tmp[9610]*kernel[6]+tmp[9611]*kernel[7]+tmp[9612]*kernel[8];
				ans[9512]<=tmp[9411]*kernel[0]+tmp[9412]*kernel[1]+tmp[9413]*kernel[2]+tmp[9511]*kernel[3]+tmp[9512]*kernel[4]+tmp[9513]*kernel[5]+tmp[9611]*kernel[6]+tmp[9612]*kernel[7]+tmp[9613]*kernel[8];
				ans[9513]<=tmp[9412]*kernel[0]+tmp[9413]*kernel[1]+tmp[9414]*kernel[2]+tmp[9512]*kernel[3]+tmp[9513]*kernel[4]+tmp[9514]*kernel[5]+tmp[9612]*kernel[6]+tmp[9613]*kernel[7]+tmp[9614]*kernel[8];
				ans[9514]<=tmp[9413]*kernel[0]+tmp[9414]*kernel[1]+tmp[9415]*kernel[2]+tmp[9513]*kernel[3]+tmp[9514]*kernel[4]+tmp[9515]*kernel[5]+tmp[9613]*kernel[6]+tmp[9614]*kernel[7]+tmp[9615]*kernel[8];
				ans[9515]<=tmp[9414]*kernel[0]+tmp[9415]*kernel[1]+tmp[9416]*kernel[2]+tmp[9514]*kernel[3]+tmp[9515]*kernel[4]+tmp[9516]*kernel[5]+tmp[9614]*kernel[6]+tmp[9615]*kernel[7]+tmp[9616]*kernel[8];
				ans[9516]<=tmp[9415]*kernel[0]+tmp[9416]*kernel[1]+tmp[9417]*kernel[2]+tmp[9515]*kernel[3]+tmp[9516]*kernel[4]+tmp[9517]*kernel[5]+tmp[9615]*kernel[6]+tmp[9616]*kernel[7]+tmp[9617]*kernel[8];
				ans[9517]<=tmp[9416]*kernel[0]+tmp[9417]*kernel[1]+tmp[9418]*kernel[2]+tmp[9516]*kernel[3]+tmp[9517]*kernel[4]+tmp[9518]*kernel[5]+tmp[9616]*kernel[6]+tmp[9617]*kernel[7]+tmp[9618]*kernel[8];
				ans[9518]<=tmp[9417]*kernel[0]+tmp[9418]*kernel[1]+tmp[9419]*kernel[2]+tmp[9517]*kernel[3]+tmp[9518]*kernel[4]+tmp[9519]*kernel[5]+tmp[9617]*kernel[6]+tmp[9618]*kernel[7]+tmp[9619]*kernel[8];
				ans[9519]<=tmp[9418]*kernel[0]+tmp[9419]*kernel[1]+tmp[9420]*kernel[2]+tmp[9518]*kernel[3]+tmp[9519]*kernel[4]+tmp[9520]*kernel[5]+tmp[9618]*kernel[6]+tmp[9619]*kernel[7]+tmp[9620]*kernel[8];
				ans[9520]<=tmp[9419]*kernel[0]+tmp[9420]*kernel[1]+tmp[9421]*kernel[2]+tmp[9519]*kernel[3]+tmp[9520]*kernel[4]+tmp[9521]*kernel[5]+tmp[9619]*kernel[6]+tmp[9620]*kernel[7]+tmp[9621]*kernel[8];
				ans[9521]<=tmp[9420]*kernel[0]+tmp[9421]*kernel[1]+tmp[9422]*kernel[2]+tmp[9520]*kernel[3]+tmp[9521]*kernel[4]+tmp[9522]*kernel[5]+tmp[9620]*kernel[6]+tmp[9621]*kernel[7]+tmp[9622]*kernel[8];
				ans[9522]<=tmp[9421]*kernel[0]+tmp[9422]*kernel[1]+tmp[9423]*kernel[2]+tmp[9521]*kernel[3]+tmp[9522]*kernel[4]+tmp[9523]*kernel[5]+tmp[9621]*kernel[6]+tmp[9622]*kernel[7]+tmp[9623]*kernel[8];
				ans[9523]<=tmp[9422]*kernel[0]+tmp[9423]*kernel[1]+tmp[9424]*kernel[2]+tmp[9522]*kernel[3]+tmp[9523]*kernel[4]+tmp[9524]*kernel[5]+tmp[9622]*kernel[6]+tmp[9623]*kernel[7]+tmp[9624]*kernel[8];
				ans[9524]<=tmp[9423]*kernel[0]+tmp[9424]*kernel[1]+tmp[9425]*kernel[2]+tmp[9523]*kernel[3]+tmp[9524]*kernel[4]+tmp[9525]*kernel[5]+tmp[9623]*kernel[6]+tmp[9624]*kernel[7]+tmp[9625]*kernel[8];
				ans[9525]<=tmp[9424]*kernel[0]+tmp[9425]*kernel[1]+tmp[9426]*kernel[2]+tmp[9524]*kernel[3]+tmp[9525]*kernel[4]+tmp[9526]*kernel[5]+tmp[9624]*kernel[6]+tmp[9625]*kernel[7]+tmp[9626]*kernel[8];
				ans[9526]<=tmp[9425]*kernel[0]+tmp[9426]*kernel[1]+tmp[9427]*kernel[2]+tmp[9525]*kernel[3]+tmp[9526]*kernel[4]+tmp[9527]*kernel[5]+tmp[9625]*kernel[6]+tmp[9626]*kernel[7]+tmp[9627]*kernel[8];
				ans[9527]<=tmp[9426]*kernel[0]+tmp[9427]*kernel[1]+tmp[9428]*kernel[2]+tmp[9526]*kernel[3]+tmp[9527]*kernel[4]+tmp[9528]*kernel[5]+tmp[9626]*kernel[6]+tmp[9627]*kernel[7]+tmp[9628]*kernel[8];
				ans[9528]<=tmp[9427]*kernel[0]+tmp[9428]*kernel[1]+tmp[9429]*kernel[2]+tmp[9527]*kernel[3]+tmp[9528]*kernel[4]+tmp[9529]*kernel[5]+tmp[9627]*kernel[6]+tmp[9628]*kernel[7]+tmp[9629]*kernel[8];
				ans[9529]<=tmp[9428]*kernel[0]+tmp[9429]*kernel[1]+tmp[9430]*kernel[2]+tmp[9528]*kernel[3]+tmp[9529]*kernel[4]+tmp[9530]*kernel[5]+tmp[9628]*kernel[6]+tmp[9629]*kernel[7]+tmp[9630]*kernel[8];
				ans[9530]<=tmp[9429]*kernel[0]+tmp[9430]*kernel[1]+tmp[9431]*kernel[2]+tmp[9529]*kernel[3]+tmp[9530]*kernel[4]+tmp[9531]*kernel[5]+tmp[9629]*kernel[6]+tmp[9630]*kernel[7]+tmp[9631]*kernel[8];
				ans[9531]<=tmp[9430]*kernel[0]+tmp[9431]*kernel[1]+tmp[9432]*kernel[2]+tmp[9530]*kernel[3]+tmp[9531]*kernel[4]+tmp[9532]*kernel[5]+tmp[9630]*kernel[6]+tmp[9631]*kernel[7]+tmp[9632]*kernel[8];
				ans[9532]<=tmp[9431]*kernel[0]+tmp[9432]*kernel[1]+tmp[9433]*kernel[2]+tmp[9531]*kernel[3]+tmp[9532]*kernel[4]+tmp[9533]*kernel[5]+tmp[9631]*kernel[6]+tmp[9632]*kernel[7]+tmp[9633]*kernel[8];
				ans[9533]<=tmp[9432]*kernel[0]+tmp[9433]*kernel[1]+tmp[9434]*kernel[2]+tmp[9532]*kernel[3]+tmp[9533]*kernel[4]+tmp[9534]*kernel[5]+tmp[9632]*kernel[6]+tmp[9633]*kernel[7]+tmp[9634]*kernel[8];
				ans[9534]<=tmp[9433]*kernel[0]+tmp[9434]*kernel[1]+tmp[9435]*kernel[2]+tmp[9533]*kernel[3]+tmp[9534]*kernel[4]+tmp[9535]*kernel[5]+tmp[9633]*kernel[6]+tmp[9634]*kernel[7]+tmp[9635]*kernel[8];
				ans[9535]<=tmp[9434]*kernel[0]+tmp[9435]*kernel[1]+tmp[9436]*kernel[2]+tmp[9534]*kernel[3]+tmp[9535]*kernel[4]+tmp[9536]*kernel[5]+tmp[9634]*kernel[6]+tmp[9635]*kernel[7]+tmp[9636]*kernel[8];
				ans[9536]<=tmp[9435]*kernel[0]+tmp[9436]*kernel[1]+tmp[9437]*kernel[2]+tmp[9535]*kernel[3]+tmp[9536]*kernel[4]+tmp[9537]*kernel[5]+tmp[9635]*kernel[6]+tmp[9636]*kernel[7]+tmp[9637]*kernel[8];
				ans[9537]<=tmp[9436]*kernel[0]+tmp[9437]*kernel[1]+tmp[9438]*kernel[2]+tmp[9536]*kernel[3]+tmp[9537]*kernel[4]+tmp[9538]*kernel[5]+tmp[9636]*kernel[6]+tmp[9637]*kernel[7]+tmp[9638]*kernel[8];
				ans[9538]<=tmp[9437]*kernel[0]+tmp[9438]*kernel[1]+tmp[9439]*kernel[2]+tmp[9537]*kernel[3]+tmp[9538]*kernel[4]+tmp[9539]*kernel[5]+tmp[9637]*kernel[6]+tmp[9638]*kernel[7]+tmp[9639]*kernel[8];
				ans[9539]<=tmp[9438]*kernel[0]+tmp[9439]*kernel[1]+tmp[9440]*kernel[2]+tmp[9538]*kernel[3]+tmp[9539]*kernel[4]+tmp[9540]*kernel[5]+tmp[9638]*kernel[6]+tmp[9639]*kernel[7]+tmp[9640]*kernel[8];
				ans[9540]<=tmp[9439]*kernel[0]+tmp[9440]*kernel[1]+tmp[9441]*kernel[2]+tmp[9539]*kernel[3]+tmp[9540]*kernel[4]+tmp[9541]*kernel[5]+tmp[9639]*kernel[6]+tmp[9640]*kernel[7]+tmp[9641]*kernel[8];
				ans[9541]<=tmp[9440]*kernel[0]+tmp[9441]*kernel[1]+tmp[9442]*kernel[2]+tmp[9540]*kernel[3]+tmp[9541]*kernel[4]+tmp[9542]*kernel[5]+tmp[9640]*kernel[6]+tmp[9641]*kernel[7]+tmp[9642]*kernel[8];
				ans[9542]<=tmp[9441]*kernel[0]+tmp[9442]*kernel[1]+tmp[9443]*kernel[2]+tmp[9541]*kernel[3]+tmp[9542]*kernel[4]+tmp[9543]*kernel[5]+tmp[9641]*kernel[6]+tmp[9642]*kernel[7]+tmp[9643]*kernel[8];
				ans[9543]<=tmp[9442]*kernel[0]+tmp[9443]*kernel[1]+tmp[9444]*kernel[2]+tmp[9542]*kernel[3]+tmp[9543]*kernel[4]+tmp[9544]*kernel[5]+tmp[9642]*kernel[6]+tmp[9643]*kernel[7]+tmp[9644]*kernel[8];
				ans[9544]<=tmp[9443]*kernel[0]+tmp[9444]*kernel[1]+tmp[9445]*kernel[2]+tmp[9543]*kernel[3]+tmp[9544]*kernel[4]+tmp[9545]*kernel[5]+tmp[9643]*kernel[6]+tmp[9644]*kernel[7]+tmp[9645]*kernel[8];
				ans[9545]<=tmp[9444]*kernel[0]+tmp[9445]*kernel[1]+tmp[9446]*kernel[2]+tmp[9544]*kernel[3]+tmp[9545]*kernel[4]+tmp[9546]*kernel[5]+tmp[9644]*kernel[6]+tmp[9645]*kernel[7]+tmp[9646]*kernel[8];
				ans[9546]<=tmp[9445]*kernel[0]+tmp[9446]*kernel[1]+tmp[9447]*kernel[2]+tmp[9545]*kernel[3]+tmp[9546]*kernel[4]+tmp[9547]*kernel[5]+tmp[9645]*kernel[6]+tmp[9646]*kernel[7]+tmp[9647]*kernel[8];
				ans[9547]<=tmp[9446]*kernel[0]+tmp[9447]*kernel[1]+tmp[9448]*kernel[2]+tmp[9546]*kernel[3]+tmp[9547]*kernel[4]+tmp[9548]*kernel[5]+tmp[9646]*kernel[6]+tmp[9647]*kernel[7]+tmp[9648]*kernel[8];
				ans[9548]<=tmp[9447]*kernel[0]+tmp[9448]*kernel[1]+tmp[9449]*kernel[2]+tmp[9547]*kernel[3]+tmp[9548]*kernel[4]+tmp[9549]*kernel[5]+tmp[9647]*kernel[6]+tmp[9648]*kernel[7]+tmp[9649]*kernel[8];
				ans[9549]<=tmp[9448]*kernel[0]+tmp[9449]*kernel[1]+tmp[9450]*kernel[2]+tmp[9548]*kernel[3]+tmp[9549]*kernel[4]+tmp[9550]*kernel[5]+tmp[9648]*kernel[6]+tmp[9649]*kernel[7]+tmp[9650]*kernel[8];
				ans[9550]<=tmp[9449]*kernel[0]+tmp[9450]*kernel[1]+tmp[9451]*kernel[2]+tmp[9549]*kernel[3]+tmp[9550]*kernel[4]+tmp[9551]*kernel[5]+tmp[9649]*kernel[6]+tmp[9650]*kernel[7]+tmp[9651]*kernel[8];
				ans[9551]<=tmp[9450]*kernel[0]+tmp[9451]*kernel[1]+tmp[9452]*kernel[2]+tmp[9550]*kernel[3]+tmp[9551]*kernel[4]+tmp[9552]*kernel[5]+tmp[9650]*kernel[6]+tmp[9651]*kernel[7]+tmp[9652]*kernel[8];
				ans[9552]<=tmp[9451]*kernel[0]+tmp[9452]*kernel[1]+tmp[9453]*kernel[2]+tmp[9551]*kernel[3]+tmp[9552]*kernel[4]+tmp[9553]*kernel[5]+tmp[9651]*kernel[6]+tmp[9652]*kernel[7]+tmp[9653]*kernel[8];
				ans[9553]<=tmp[9452]*kernel[0]+tmp[9453]*kernel[1]+tmp[9454]*kernel[2]+tmp[9552]*kernel[3]+tmp[9553]*kernel[4]+tmp[9554]*kernel[5]+tmp[9652]*kernel[6]+tmp[9653]*kernel[7]+tmp[9654]*kernel[8];
				ans[9554]<=tmp[9453]*kernel[0]+tmp[9454]*kernel[1]+tmp[9455]*kernel[2]+tmp[9553]*kernel[3]+tmp[9554]*kernel[4]+tmp[9555]*kernel[5]+tmp[9653]*kernel[6]+tmp[9654]*kernel[7]+tmp[9655]*kernel[8];
				ans[9555]<=tmp[9454]*kernel[0]+tmp[9455]*kernel[1]+tmp[9456]*kernel[2]+tmp[9554]*kernel[3]+tmp[9555]*kernel[4]+tmp[9556]*kernel[5]+tmp[9654]*kernel[6]+tmp[9655]*kernel[7]+tmp[9656]*kernel[8];
				ans[9556]<=tmp[9455]*kernel[0]+tmp[9456]*kernel[1]+tmp[9457]*kernel[2]+tmp[9555]*kernel[3]+tmp[9556]*kernel[4]+tmp[9557]*kernel[5]+tmp[9655]*kernel[6]+tmp[9656]*kernel[7]+tmp[9657]*kernel[8];
				ans[9557]<=tmp[9456]*kernel[0]+tmp[9457]*kernel[1]+tmp[9458]*kernel[2]+tmp[9556]*kernel[3]+tmp[9557]*kernel[4]+tmp[9558]*kernel[5]+tmp[9656]*kernel[6]+tmp[9657]*kernel[7]+tmp[9658]*kernel[8];
				ans[9558]<=tmp[9457]*kernel[0]+tmp[9458]*kernel[1]+tmp[9459]*kernel[2]+tmp[9557]*kernel[3]+tmp[9558]*kernel[4]+tmp[9559]*kernel[5]+tmp[9657]*kernel[6]+tmp[9658]*kernel[7]+tmp[9659]*kernel[8];
				ans[9559]<=tmp[9458]*kernel[0]+tmp[9459]*kernel[1]+tmp[9460]*kernel[2]+tmp[9558]*kernel[3]+tmp[9559]*kernel[4]+tmp[9560]*kernel[5]+tmp[9658]*kernel[6]+tmp[9659]*kernel[7]+tmp[9660]*kernel[8];
				ans[9560]<=tmp[9459]*kernel[0]+tmp[9460]*kernel[1]+tmp[9461]*kernel[2]+tmp[9559]*kernel[3]+tmp[9560]*kernel[4]+tmp[9561]*kernel[5]+tmp[9659]*kernel[6]+tmp[9660]*kernel[7]+tmp[9661]*kernel[8];
				ans[9561]<=tmp[9460]*kernel[0]+tmp[9461]*kernel[1]+tmp[9462]*kernel[2]+tmp[9560]*kernel[3]+tmp[9561]*kernel[4]+tmp[9562]*kernel[5]+tmp[9660]*kernel[6]+tmp[9661]*kernel[7]+tmp[9662]*kernel[8];
				ans[9562]<=tmp[9461]*kernel[0]+tmp[9462]*kernel[1]+tmp[9463]*kernel[2]+tmp[9561]*kernel[3]+tmp[9562]*kernel[4]+tmp[9563]*kernel[5]+tmp[9661]*kernel[6]+tmp[9662]*kernel[7]+tmp[9663]*kernel[8];
				ans[9563]<=tmp[9462]*kernel[0]+tmp[9463]*kernel[1]+tmp[9464]*kernel[2]+tmp[9562]*kernel[3]+tmp[9563]*kernel[4]+tmp[9564]*kernel[5]+tmp[9662]*kernel[6]+tmp[9663]*kernel[7]+tmp[9664]*kernel[8];
				ans[9564]<=tmp[9463]*kernel[0]+tmp[9464]*kernel[1]+tmp[9465]*kernel[2]+tmp[9563]*kernel[3]+tmp[9564]*kernel[4]+tmp[9565]*kernel[5]+tmp[9663]*kernel[6]+tmp[9664]*kernel[7]+tmp[9665]*kernel[8];
				ans[9565]<=tmp[9464]*kernel[0]+tmp[9465]*kernel[1]+tmp[9466]*kernel[2]+tmp[9564]*kernel[3]+tmp[9565]*kernel[4]+tmp[9566]*kernel[5]+tmp[9664]*kernel[6]+tmp[9665]*kernel[7]+tmp[9666]*kernel[8];
				ans[9566]<=tmp[9465]*kernel[0]+tmp[9466]*kernel[1]+tmp[9467]*kernel[2]+tmp[9565]*kernel[3]+tmp[9566]*kernel[4]+tmp[9567]*kernel[5]+tmp[9665]*kernel[6]+tmp[9666]*kernel[7]+tmp[9667]*kernel[8];
				ans[9567]<=tmp[9466]*kernel[0]+tmp[9467]*kernel[1]+tmp[9468]*kernel[2]+tmp[9566]*kernel[3]+tmp[9567]*kernel[4]+tmp[9568]*kernel[5]+tmp[9666]*kernel[6]+tmp[9667]*kernel[7]+tmp[9668]*kernel[8];
				ans[9568]<=tmp[9467]*kernel[0]+tmp[9468]*kernel[1]+tmp[9469]*kernel[2]+tmp[9567]*kernel[3]+tmp[9568]*kernel[4]+tmp[9569]*kernel[5]+tmp[9667]*kernel[6]+tmp[9668]*kernel[7]+tmp[9669]*kernel[8];
				ans[9569]<=tmp[9468]*kernel[0]+tmp[9469]*kernel[1]+tmp[9470]*kernel[2]+tmp[9568]*kernel[3]+tmp[9569]*kernel[4]+tmp[9570]*kernel[5]+tmp[9668]*kernel[6]+tmp[9669]*kernel[7]+tmp[9670]*kernel[8];
				ans[9570]<=tmp[9469]*kernel[0]+tmp[9470]*kernel[1]+tmp[9471]*kernel[2]+tmp[9569]*kernel[3]+tmp[9570]*kernel[4]+tmp[9571]*kernel[5]+tmp[9669]*kernel[6]+tmp[9670]*kernel[7]+tmp[9671]*kernel[8];
				ans[9571]<=tmp[9470]*kernel[0]+tmp[9471]*kernel[1]+tmp[9472]*kernel[2]+tmp[9570]*kernel[3]+tmp[9571]*kernel[4]+tmp[9572]*kernel[5]+tmp[9670]*kernel[6]+tmp[9671]*kernel[7]+tmp[9672]*kernel[8];
				ans[9572]<=tmp[9471]*kernel[0]+tmp[9472]*kernel[1]+tmp[9473]*kernel[2]+tmp[9571]*kernel[3]+tmp[9572]*kernel[4]+tmp[9573]*kernel[5]+tmp[9671]*kernel[6]+tmp[9672]*kernel[7]+tmp[9673]*kernel[8];
				ans[9573]<=tmp[9472]*kernel[0]+tmp[9473]*kernel[1]+tmp[9474]*kernel[2]+tmp[9572]*kernel[3]+tmp[9573]*kernel[4]+tmp[9574]*kernel[5]+tmp[9672]*kernel[6]+tmp[9673]*kernel[7]+tmp[9674]*kernel[8];
				ans[9574]<=tmp[9473]*kernel[0]+tmp[9474]*kernel[1]+tmp[9475]*kernel[2]+tmp[9573]*kernel[3]+tmp[9574]*kernel[4]+tmp[9575]*kernel[5]+tmp[9673]*kernel[6]+tmp[9674]*kernel[7]+tmp[9675]*kernel[8];
				ans[9575]<=tmp[9474]*kernel[0]+tmp[9475]*kernel[1]+tmp[9476]*kernel[2]+tmp[9574]*kernel[3]+tmp[9575]*kernel[4]+tmp[9576]*kernel[5]+tmp[9674]*kernel[6]+tmp[9675]*kernel[7]+tmp[9676]*kernel[8];
				ans[9576]<=tmp[9475]*kernel[0]+tmp[9476]*kernel[1]+tmp[9477]*kernel[2]+tmp[9575]*kernel[3]+tmp[9576]*kernel[4]+tmp[9577]*kernel[5]+tmp[9675]*kernel[6]+tmp[9676]*kernel[7]+tmp[9677]*kernel[8];
				ans[9577]<=tmp[9476]*kernel[0]+tmp[9477]*kernel[1]+tmp[9478]*kernel[2]+tmp[9576]*kernel[3]+tmp[9577]*kernel[4]+tmp[9578]*kernel[5]+tmp[9676]*kernel[6]+tmp[9677]*kernel[7]+tmp[9678]*kernel[8];
				ans[9578]<=tmp[9477]*kernel[0]+tmp[9478]*kernel[1]+tmp[9479]*kernel[2]+tmp[9577]*kernel[3]+tmp[9578]*kernel[4]+tmp[9579]*kernel[5]+tmp[9677]*kernel[6]+tmp[9678]*kernel[7]+tmp[9679]*kernel[8];
				ans[9579]<=tmp[9478]*kernel[0]+tmp[9479]*kernel[1]+tmp[9480]*kernel[2]+tmp[9578]*kernel[3]+tmp[9579]*kernel[4]+tmp[9580]*kernel[5]+tmp[9678]*kernel[6]+tmp[9679]*kernel[7]+tmp[9680]*kernel[8];
				ans[9580]<=tmp[9479]*kernel[0]+tmp[9480]*kernel[1]+tmp[9481]*kernel[2]+tmp[9579]*kernel[3]+tmp[9580]*kernel[4]+tmp[9581]*kernel[5]+tmp[9679]*kernel[6]+tmp[9680]*kernel[7]+tmp[9681]*kernel[8];
				ans[9581]<=tmp[9480]*kernel[0]+tmp[9481]*kernel[1]+tmp[9482]*kernel[2]+tmp[9580]*kernel[3]+tmp[9581]*kernel[4]+tmp[9582]*kernel[5]+tmp[9680]*kernel[6]+tmp[9681]*kernel[7]+tmp[9682]*kernel[8];
				ans[9582]<=tmp[9481]*kernel[0]+tmp[9482]*kernel[1]+tmp[9483]*kernel[2]+tmp[9581]*kernel[3]+tmp[9582]*kernel[4]+tmp[9583]*kernel[5]+tmp[9681]*kernel[6]+tmp[9682]*kernel[7]+tmp[9683]*kernel[8];
				ans[9583]<=tmp[9482]*kernel[0]+tmp[9483]*kernel[1]+tmp[9484]*kernel[2]+tmp[9582]*kernel[3]+tmp[9583]*kernel[4]+tmp[9584]*kernel[5]+tmp[9682]*kernel[6]+tmp[9683]*kernel[7]+tmp[9684]*kernel[8];
				ans[9584]<=tmp[9483]*kernel[0]+tmp[9484]*kernel[1]+tmp[9485]*kernel[2]+tmp[9583]*kernel[3]+tmp[9584]*kernel[4]+tmp[9585]*kernel[5]+tmp[9683]*kernel[6]+tmp[9684]*kernel[7]+tmp[9685]*kernel[8];
				ans[9585]<=tmp[9484]*kernel[0]+tmp[9485]*kernel[1]+tmp[9486]*kernel[2]+tmp[9584]*kernel[3]+tmp[9585]*kernel[4]+tmp[9586]*kernel[5]+tmp[9684]*kernel[6]+tmp[9685]*kernel[7]+tmp[9686]*kernel[8];
				ans[9586]<=tmp[9485]*kernel[0]+tmp[9486]*kernel[1]+tmp[9487]*kernel[2]+tmp[9585]*kernel[3]+tmp[9586]*kernel[4]+tmp[9587]*kernel[5]+tmp[9685]*kernel[6]+tmp[9686]*kernel[7]+tmp[9687]*kernel[8];
				ans[9587]<=tmp[9486]*kernel[0]+tmp[9487]*kernel[1]+tmp[9488]*kernel[2]+tmp[9586]*kernel[3]+tmp[9587]*kernel[4]+tmp[9588]*kernel[5]+tmp[9686]*kernel[6]+tmp[9687]*kernel[7]+tmp[9688]*kernel[8];
				ans[9588]<=tmp[9487]*kernel[0]+tmp[9488]*kernel[1]+tmp[9489]*kernel[2]+tmp[9587]*kernel[3]+tmp[9588]*kernel[4]+tmp[9589]*kernel[5]+tmp[9687]*kernel[6]+tmp[9688]*kernel[7]+tmp[9689]*kernel[8];
				ans[9589]<=tmp[9488]*kernel[0]+tmp[9489]*kernel[1]+tmp[9490]*kernel[2]+tmp[9588]*kernel[3]+tmp[9589]*kernel[4]+tmp[9590]*kernel[5]+tmp[9688]*kernel[6]+tmp[9689]*kernel[7]+tmp[9690]*kernel[8];
				ans[9590]<=tmp[9489]*kernel[0]+tmp[9490]*kernel[1]+tmp[9491]*kernel[2]+tmp[9589]*kernel[3]+tmp[9590]*kernel[4]+tmp[9591]*kernel[5]+tmp[9689]*kernel[6]+tmp[9690]*kernel[7]+tmp[9691]*kernel[8];
				ans[9591]<=tmp[9490]*kernel[0]+tmp[9491]*kernel[1]+tmp[9492]*kernel[2]+tmp[9590]*kernel[3]+tmp[9591]*kernel[4]+tmp[9592]*kernel[5]+tmp[9690]*kernel[6]+tmp[9691]*kernel[7]+tmp[9692]*kernel[8];
				ans[9592]<=tmp[9491]*kernel[0]+tmp[9492]*kernel[1]+tmp[9493]*kernel[2]+tmp[9591]*kernel[3]+tmp[9592]*kernel[4]+tmp[9593]*kernel[5]+tmp[9691]*kernel[6]+tmp[9692]*kernel[7]+tmp[9693]*kernel[8];
				ans[9593]<=tmp[9492]*kernel[0]+tmp[9493]*kernel[1]+tmp[9494]*kernel[2]+tmp[9592]*kernel[3]+tmp[9593]*kernel[4]+tmp[9594]*kernel[5]+tmp[9692]*kernel[6]+tmp[9693]*kernel[7]+tmp[9694]*kernel[8];
				ans[9594]<=tmp[9493]*kernel[0]+tmp[9494]*kernel[1]+tmp[9495]*kernel[2]+tmp[9593]*kernel[3]+tmp[9594]*kernel[4]+tmp[9595]*kernel[5]+tmp[9693]*kernel[6]+tmp[9694]*kernel[7]+tmp[9695]*kernel[8];
				ans[9595]<=tmp[9494]*kernel[0]+tmp[9495]*kernel[1]+tmp[9496]*kernel[2]+tmp[9594]*kernel[3]+tmp[9595]*kernel[4]+tmp[9596]*kernel[5]+tmp[9694]*kernel[6]+tmp[9695]*kernel[7]+tmp[9696]*kernel[8];
				ans[9596]<=tmp[9495]*kernel[0]+tmp[9496]*kernel[1]+tmp[9497]*kernel[2]+tmp[9595]*kernel[3]+tmp[9596]*kernel[4]+tmp[9597]*kernel[5]+tmp[9695]*kernel[6]+tmp[9696]*kernel[7]+tmp[9697]*kernel[8];
				ans[9597]<=tmp[9496]*kernel[0]+tmp[9497]*kernel[1]+tmp[9498]*kernel[2]+tmp[9596]*kernel[3]+tmp[9597]*kernel[4]+tmp[9598]*kernel[5]+tmp[9696]*kernel[6]+tmp[9697]*kernel[7]+tmp[9698]*kernel[8];
				ans[9598]<=tmp[9497]*kernel[0]+tmp[9498]*kernel[1]+tmp[9499]*kernel[2]+tmp[9597]*kernel[3]+tmp[9598]*kernel[4]+tmp[9599]*kernel[5]+tmp[9697]*kernel[6]+tmp[9698]*kernel[7]+tmp[9699]*kernel[8];
				ans[9599]<=tmp[9498]*kernel[0]+tmp[9499]*kernel[1]+tmp[9598]*kernel[3]+tmp[9599]*kernel[4]+tmp[9698]*kernel[6]+tmp[9699]*kernel[7];
				ans[9600]<=tmp[9500]*kernel[1]+tmp[9501]*kernel[2]+tmp[9600]*kernel[4]+tmp[9601]*kernel[5]+tmp[9700]*kernel[7]+tmp[9701]*kernel[8];
				ans[9601]<=tmp[9500]*kernel[0]+tmp[9501]*kernel[1]+tmp[9502]*kernel[2]+tmp[9600]*kernel[3]+tmp[9601]*kernel[4]+tmp[9602]*kernel[5]+tmp[9700]*kernel[6]+tmp[9701]*kernel[7]+tmp[9702]*kernel[8];
				ans[9602]<=tmp[9501]*kernel[0]+tmp[9502]*kernel[1]+tmp[9503]*kernel[2]+tmp[9601]*kernel[3]+tmp[9602]*kernel[4]+tmp[9603]*kernel[5]+tmp[9701]*kernel[6]+tmp[9702]*kernel[7]+tmp[9703]*kernel[8];
				ans[9603]<=tmp[9502]*kernel[0]+tmp[9503]*kernel[1]+tmp[9504]*kernel[2]+tmp[9602]*kernel[3]+tmp[9603]*kernel[4]+tmp[9604]*kernel[5]+tmp[9702]*kernel[6]+tmp[9703]*kernel[7]+tmp[9704]*kernel[8];
				ans[9604]<=tmp[9503]*kernel[0]+tmp[9504]*kernel[1]+tmp[9505]*kernel[2]+tmp[9603]*kernel[3]+tmp[9604]*kernel[4]+tmp[9605]*kernel[5]+tmp[9703]*kernel[6]+tmp[9704]*kernel[7]+tmp[9705]*kernel[8];
				ans[9605]<=tmp[9504]*kernel[0]+tmp[9505]*kernel[1]+tmp[9506]*kernel[2]+tmp[9604]*kernel[3]+tmp[9605]*kernel[4]+tmp[9606]*kernel[5]+tmp[9704]*kernel[6]+tmp[9705]*kernel[7]+tmp[9706]*kernel[8];
				ans[9606]<=tmp[9505]*kernel[0]+tmp[9506]*kernel[1]+tmp[9507]*kernel[2]+tmp[9605]*kernel[3]+tmp[9606]*kernel[4]+tmp[9607]*kernel[5]+tmp[9705]*kernel[6]+tmp[9706]*kernel[7]+tmp[9707]*kernel[8];
				ans[9607]<=tmp[9506]*kernel[0]+tmp[9507]*kernel[1]+tmp[9508]*kernel[2]+tmp[9606]*kernel[3]+tmp[9607]*kernel[4]+tmp[9608]*kernel[5]+tmp[9706]*kernel[6]+tmp[9707]*kernel[7]+tmp[9708]*kernel[8];
				ans[9608]<=tmp[9507]*kernel[0]+tmp[9508]*kernel[1]+tmp[9509]*kernel[2]+tmp[9607]*kernel[3]+tmp[9608]*kernel[4]+tmp[9609]*kernel[5]+tmp[9707]*kernel[6]+tmp[9708]*kernel[7]+tmp[9709]*kernel[8];
				ans[9609]<=tmp[9508]*kernel[0]+tmp[9509]*kernel[1]+tmp[9510]*kernel[2]+tmp[9608]*kernel[3]+tmp[9609]*kernel[4]+tmp[9610]*kernel[5]+tmp[9708]*kernel[6]+tmp[9709]*kernel[7]+tmp[9710]*kernel[8];
				ans[9610]<=tmp[9509]*kernel[0]+tmp[9510]*kernel[1]+tmp[9511]*kernel[2]+tmp[9609]*kernel[3]+tmp[9610]*kernel[4]+tmp[9611]*kernel[5]+tmp[9709]*kernel[6]+tmp[9710]*kernel[7]+tmp[9711]*kernel[8];
				ans[9611]<=tmp[9510]*kernel[0]+tmp[9511]*kernel[1]+tmp[9512]*kernel[2]+tmp[9610]*kernel[3]+tmp[9611]*kernel[4]+tmp[9612]*kernel[5]+tmp[9710]*kernel[6]+tmp[9711]*kernel[7]+tmp[9712]*kernel[8];
				ans[9612]<=tmp[9511]*kernel[0]+tmp[9512]*kernel[1]+tmp[9513]*kernel[2]+tmp[9611]*kernel[3]+tmp[9612]*kernel[4]+tmp[9613]*kernel[5]+tmp[9711]*kernel[6]+tmp[9712]*kernel[7]+tmp[9713]*kernel[8];
				ans[9613]<=tmp[9512]*kernel[0]+tmp[9513]*kernel[1]+tmp[9514]*kernel[2]+tmp[9612]*kernel[3]+tmp[9613]*kernel[4]+tmp[9614]*kernel[5]+tmp[9712]*kernel[6]+tmp[9713]*kernel[7]+tmp[9714]*kernel[8];
				ans[9614]<=tmp[9513]*kernel[0]+tmp[9514]*kernel[1]+tmp[9515]*kernel[2]+tmp[9613]*kernel[3]+tmp[9614]*kernel[4]+tmp[9615]*kernel[5]+tmp[9713]*kernel[6]+tmp[9714]*kernel[7]+tmp[9715]*kernel[8];
				ans[9615]<=tmp[9514]*kernel[0]+tmp[9515]*kernel[1]+tmp[9516]*kernel[2]+tmp[9614]*kernel[3]+tmp[9615]*kernel[4]+tmp[9616]*kernel[5]+tmp[9714]*kernel[6]+tmp[9715]*kernel[7]+tmp[9716]*kernel[8];
				ans[9616]<=tmp[9515]*kernel[0]+tmp[9516]*kernel[1]+tmp[9517]*kernel[2]+tmp[9615]*kernel[3]+tmp[9616]*kernel[4]+tmp[9617]*kernel[5]+tmp[9715]*kernel[6]+tmp[9716]*kernel[7]+tmp[9717]*kernel[8];
				ans[9617]<=tmp[9516]*kernel[0]+tmp[9517]*kernel[1]+tmp[9518]*kernel[2]+tmp[9616]*kernel[3]+tmp[9617]*kernel[4]+tmp[9618]*kernel[5]+tmp[9716]*kernel[6]+tmp[9717]*kernel[7]+tmp[9718]*kernel[8];
				ans[9618]<=tmp[9517]*kernel[0]+tmp[9518]*kernel[1]+tmp[9519]*kernel[2]+tmp[9617]*kernel[3]+tmp[9618]*kernel[4]+tmp[9619]*kernel[5]+tmp[9717]*kernel[6]+tmp[9718]*kernel[7]+tmp[9719]*kernel[8];
				ans[9619]<=tmp[9518]*kernel[0]+tmp[9519]*kernel[1]+tmp[9520]*kernel[2]+tmp[9618]*kernel[3]+tmp[9619]*kernel[4]+tmp[9620]*kernel[5]+tmp[9718]*kernel[6]+tmp[9719]*kernel[7]+tmp[9720]*kernel[8];
				ans[9620]<=tmp[9519]*kernel[0]+tmp[9520]*kernel[1]+tmp[9521]*kernel[2]+tmp[9619]*kernel[3]+tmp[9620]*kernel[4]+tmp[9621]*kernel[5]+tmp[9719]*kernel[6]+tmp[9720]*kernel[7]+tmp[9721]*kernel[8];
				ans[9621]<=tmp[9520]*kernel[0]+tmp[9521]*kernel[1]+tmp[9522]*kernel[2]+tmp[9620]*kernel[3]+tmp[9621]*kernel[4]+tmp[9622]*kernel[5]+tmp[9720]*kernel[6]+tmp[9721]*kernel[7]+tmp[9722]*kernel[8];
				ans[9622]<=tmp[9521]*kernel[0]+tmp[9522]*kernel[1]+tmp[9523]*kernel[2]+tmp[9621]*kernel[3]+tmp[9622]*kernel[4]+tmp[9623]*kernel[5]+tmp[9721]*kernel[6]+tmp[9722]*kernel[7]+tmp[9723]*kernel[8];
				ans[9623]<=tmp[9522]*kernel[0]+tmp[9523]*kernel[1]+tmp[9524]*kernel[2]+tmp[9622]*kernel[3]+tmp[9623]*kernel[4]+tmp[9624]*kernel[5]+tmp[9722]*kernel[6]+tmp[9723]*kernel[7]+tmp[9724]*kernel[8];
				ans[9624]<=tmp[9523]*kernel[0]+tmp[9524]*kernel[1]+tmp[9525]*kernel[2]+tmp[9623]*kernel[3]+tmp[9624]*kernel[4]+tmp[9625]*kernel[5]+tmp[9723]*kernel[6]+tmp[9724]*kernel[7]+tmp[9725]*kernel[8];
				ans[9625]<=tmp[9524]*kernel[0]+tmp[9525]*kernel[1]+tmp[9526]*kernel[2]+tmp[9624]*kernel[3]+tmp[9625]*kernel[4]+tmp[9626]*kernel[5]+tmp[9724]*kernel[6]+tmp[9725]*kernel[7]+tmp[9726]*kernel[8];
				ans[9626]<=tmp[9525]*kernel[0]+tmp[9526]*kernel[1]+tmp[9527]*kernel[2]+tmp[9625]*kernel[3]+tmp[9626]*kernel[4]+tmp[9627]*kernel[5]+tmp[9725]*kernel[6]+tmp[9726]*kernel[7]+tmp[9727]*kernel[8];
				ans[9627]<=tmp[9526]*kernel[0]+tmp[9527]*kernel[1]+tmp[9528]*kernel[2]+tmp[9626]*kernel[3]+tmp[9627]*kernel[4]+tmp[9628]*kernel[5]+tmp[9726]*kernel[6]+tmp[9727]*kernel[7]+tmp[9728]*kernel[8];
				ans[9628]<=tmp[9527]*kernel[0]+tmp[9528]*kernel[1]+tmp[9529]*kernel[2]+tmp[9627]*kernel[3]+tmp[9628]*kernel[4]+tmp[9629]*kernel[5]+tmp[9727]*kernel[6]+tmp[9728]*kernel[7]+tmp[9729]*kernel[8];
				ans[9629]<=tmp[9528]*kernel[0]+tmp[9529]*kernel[1]+tmp[9530]*kernel[2]+tmp[9628]*kernel[3]+tmp[9629]*kernel[4]+tmp[9630]*kernel[5]+tmp[9728]*kernel[6]+tmp[9729]*kernel[7]+tmp[9730]*kernel[8];
				ans[9630]<=tmp[9529]*kernel[0]+tmp[9530]*kernel[1]+tmp[9531]*kernel[2]+tmp[9629]*kernel[3]+tmp[9630]*kernel[4]+tmp[9631]*kernel[5]+tmp[9729]*kernel[6]+tmp[9730]*kernel[7]+tmp[9731]*kernel[8];
				ans[9631]<=tmp[9530]*kernel[0]+tmp[9531]*kernel[1]+tmp[9532]*kernel[2]+tmp[9630]*kernel[3]+tmp[9631]*kernel[4]+tmp[9632]*kernel[5]+tmp[9730]*kernel[6]+tmp[9731]*kernel[7]+tmp[9732]*kernel[8];
				ans[9632]<=tmp[9531]*kernel[0]+tmp[9532]*kernel[1]+tmp[9533]*kernel[2]+tmp[9631]*kernel[3]+tmp[9632]*kernel[4]+tmp[9633]*kernel[5]+tmp[9731]*kernel[6]+tmp[9732]*kernel[7]+tmp[9733]*kernel[8];
				ans[9633]<=tmp[9532]*kernel[0]+tmp[9533]*kernel[1]+tmp[9534]*kernel[2]+tmp[9632]*kernel[3]+tmp[9633]*kernel[4]+tmp[9634]*kernel[5]+tmp[9732]*kernel[6]+tmp[9733]*kernel[7]+tmp[9734]*kernel[8];
				ans[9634]<=tmp[9533]*kernel[0]+tmp[9534]*kernel[1]+tmp[9535]*kernel[2]+tmp[9633]*kernel[3]+tmp[9634]*kernel[4]+tmp[9635]*kernel[5]+tmp[9733]*kernel[6]+tmp[9734]*kernel[7]+tmp[9735]*kernel[8];
				ans[9635]<=tmp[9534]*kernel[0]+tmp[9535]*kernel[1]+tmp[9536]*kernel[2]+tmp[9634]*kernel[3]+tmp[9635]*kernel[4]+tmp[9636]*kernel[5]+tmp[9734]*kernel[6]+tmp[9735]*kernel[7]+tmp[9736]*kernel[8];
				ans[9636]<=tmp[9535]*kernel[0]+tmp[9536]*kernel[1]+tmp[9537]*kernel[2]+tmp[9635]*kernel[3]+tmp[9636]*kernel[4]+tmp[9637]*kernel[5]+tmp[9735]*kernel[6]+tmp[9736]*kernel[7]+tmp[9737]*kernel[8];
				ans[9637]<=tmp[9536]*kernel[0]+tmp[9537]*kernel[1]+tmp[9538]*kernel[2]+tmp[9636]*kernel[3]+tmp[9637]*kernel[4]+tmp[9638]*kernel[5]+tmp[9736]*kernel[6]+tmp[9737]*kernel[7]+tmp[9738]*kernel[8];
				ans[9638]<=tmp[9537]*kernel[0]+tmp[9538]*kernel[1]+tmp[9539]*kernel[2]+tmp[9637]*kernel[3]+tmp[9638]*kernel[4]+tmp[9639]*kernel[5]+tmp[9737]*kernel[6]+tmp[9738]*kernel[7]+tmp[9739]*kernel[8];
				ans[9639]<=tmp[9538]*kernel[0]+tmp[9539]*kernel[1]+tmp[9540]*kernel[2]+tmp[9638]*kernel[3]+tmp[9639]*kernel[4]+tmp[9640]*kernel[5]+tmp[9738]*kernel[6]+tmp[9739]*kernel[7]+tmp[9740]*kernel[8];
				ans[9640]<=tmp[9539]*kernel[0]+tmp[9540]*kernel[1]+tmp[9541]*kernel[2]+tmp[9639]*kernel[3]+tmp[9640]*kernel[4]+tmp[9641]*kernel[5]+tmp[9739]*kernel[6]+tmp[9740]*kernel[7]+tmp[9741]*kernel[8];
				ans[9641]<=tmp[9540]*kernel[0]+tmp[9541]*kernel[1]+tmp[9542]*kernel[2]+tmp[9640]*kernel[3]+tmp[9641]*kernel[4]+tmp[9642]*kernel[5]+tmp[9740]*kernel[6]+tmp[9741]*kernel[7]+tmp[9742]*kernel[8];
				ans[9642]<=tmp[9541]*kernel[0]+tmp[9542]*kernel[1]+tmp[9543]*kernel[2]+tmp[9641]*kernel[3]+tmp[9642]*kernel[4]+tmp[9643]*kernel[5]+tmp[9741]*kernel[6]+tmp[9742]*kernel[7]+tmp[9743]*kernel[8];
				ans[9643]<=tmp[9542]*kernel[0]+tmp[9543]*kernel[1]+tmp[9544]*kernel[2]+tmp[9642]*kernel[3]+tmp[9643]*kernel[4]+tmp[9644]*kernel[5]+tmp[9742]*kernel[6]+tmp[9743]*kernel[7]+tmp[9744]*kernel[8];
				ans[9644]<=tmp[9543]*kernel[0]+tmp[9544]*kernel[1]+tmp[9545]*kernel[2]+tmp[9643]*kernel[3]+tmp[9644]*kernel[4]+tmp[9645]*kernel[5]+tmp[9743]*kernel[6]+tmp[9744]*kernel[7]+tmp[9745]*kernel[8];
				ans[9645]<=tmp[9544]*kernel[0]+tmp[9545]*kernel[1]+tmp[9546]*kernel[2]+tmp[9644]*kernel[3]+tmp[9645]*kernel[4]+tmp[9646]*kernel[5]+tmp[9744]*kernel[6]+tmp[9745]*kernel[7]+tmp[9746]*kernel[8];
				ans[9646]<=tmp[9545]*kernel[0]+tmp[9546]*kernel[1]+tmp[9547]*kernel[2]+tmp[9645]*kernel[3]+tmp[9646]*kernel[4]+tmp[9647]*kernel[5]+tmp[9745]*kernel[6]+tmp[9746]*kernel[7]+tmp[9747]*kernel[8];
				ans[9647]<=tmp[9546]*kernel[0]+tmp[9547]*kernel[1]+tmp[9548]*kernel[2]+tmp[9646]*kernel[3]+tmp[9647]*kernel[4]+tmp[9648]*kernel[5]+tmp[9746]*kernel[6]+tmp[9747]*kernel[7]+tmp[9748]*kernel[8];
				ans[9648]<=tmp[9547]*kernel[0]+tmp[9548]*kernel[1]+tmp[9549]*kernel[2]+tmp[9647]*kernel[3]+tmp[9648]*kernel[4]+tmp[9649]*kernel[5]+tmp[9747]*kernel[6]+tmp[9748]*kernel[7]+tmp[9749]*kernel[8];
				ans[9649]<=tmp[9548]*kernel[0]+tmp[9549]*kernel[1]+tmp[9550]*kernel[2]+tmp[9648]*kernel[3]+tmp[9649]*kernel[4]+tmp[9650]*kernel[5]+tmp[9748]*kernel[6]+tmp[9749]*kernel[7]+tmp[9750]*kernel[8];
				ans[9650]<=tmp[9549]*kernel[0]+tmp[9550]*kernel[1]+tmp[9551]*kernel[2]+tmp[9649]*kernel[3]+tmp[9650]*kernel[4]+tmp[9651]*kernel[5]+tmp[9749]*kernel[6]+tmp[9750]*kernel[7]+tmp[9751]*kernel[8];
				ans[9651]<=tmp[9550]*kernel[0]+tmp[9551]*kernel[1]+tmp[9552]*kernel[2]+tmp[9650]*kernel[3]+tmp[9651]*kernel[4]+tmp[9652]*kernel[5]+tmp[9750]*kernel[6]+tmp[9751]*kernel[7]+tmp[9752]*kernel[8];
				ans[9652]<=tmp[9551]*kernel[0]+tmp[9552]*kernel[1]+tmp[9553]*kernel[2]+tmp[9651]*kernel[3]+tmp[9652]*kernel[4]+tmp[9653]*kernel[5]+tmp[9751]*kernel[6]+tmp[9752]*kernel[7]+tmp[9753]*kernel[8];
				ans[9653]<=tmp[9552]*kernel[0]+tmp[9553]*kernel[1]+tmp[9554]*kernel[2]+tmp[9652]*kernel[3]+tmp[9653]*kernel[4]+tmp[9654]*kernel[5]+tmp[9752]*kernel[6]+tmp[9753]*kernel[7]+tmp[9754]*kernel[8];
				ans[9654]<=tmp[9553]*kernel[0]+tmp[9554]*kernel[1]+tmp[9555]*kernel[2]+tmp[9653]*kernel[3]+tmp[9654]*kernel[4]+tmp[9655]*kernel[5]+tmp[9753]*kernel[6]+tmp[9754]*kernel[7]+tmp[9755]*kernel[8];
				ans[9655]<=tmp[9554]*kernel[0]+tmp[9555]*kernel[1]+tmp[9556]*kernel[2]+tmp[9654]*kernel[3]+tmp[9655]*kernel[4]+tmp[9656]*kernel[5]+tmp[9754]*kernel[6]+tmp[9755]*kernel[7]+tmp[9756]*kernel[8];
				ans[9656]<=tmp[9555]*kernel[0]+tmp[9556]*kernel[1]+tmp[9557]*kernel[2]+tmp[9655]*kernel[3]+tmp[9656]*kernel[4]+tmp[9657]*kernel[5]+tmp[9755]*kernel[6]+tmp[9756]*kernel[7]+tmp[9757]*kernel[8];
				ans[9657]<=tmp[9556]*kernel[0]+tmp[9557]*kernel[1]+tmp[9558]*kernel[2]+tmp[9656]*kernel[3]+tmp[9657]*kernel[4]+tmp[9658]*kernel[5]+tmp[9756]*kernel[6]+tmp[9757]*kernel[7]+tmp[9758]*kernel[8];
				ans[9658]<=tmp[9557]*kernel[0]+tmp[9558]*kernel[1]+tmp[9559]*kernel[2]+tmp[9657]*kernel[3]+tmp[9658]*kernel[4]+tmp[9659]*kernel[5]+tmp[9757]*kernel[6]+tmp[9758]*kernel[7]+tmp[9759]*kernel[8];
				ans[9659]<=tmp[9558]*kernel[0]+tmp[9559]*kernel[1]+tmp[9560]*kernel[2]+tmp[9658]*kernel[3]+tmp[9659]*kernel[4]+tmp[9660]*kernel[5]+tmp[9758]*kernel[6]+tmp[9759]*kernel[7]+tmp[9760]*kernel[8];
				ans[9660]<=tmp[9559]*kernel[0]+tmp[9560]*kernel[1]+tmp[9561]*kernel[2]+tmp[9659]*kernel[3]+tmp[9660]*kernel[4]+tmp[9661]*kernel[5]+tmp[9759]*kernel[6]+tmp[9760]*kernel[7]+tmp[9761]*kernel[8];
				ans[9661]<=tmp[9560]*kernel[0]+tmp[9561]*kernel[1]+tmp[9562]*kernel[2]+tmp[9660]*kernel[3]+tmp[9661]*kernel[4]+tmp[9662]*kernel[5]+tmp[9760]*kernel[6]+tmp[9761]*kernel[7]+tmp[9762]*kernel[8];
				ans[9662]<=tmp[9561]*kernel[0]+tmp[9562]*kernel[1]+tmp[9563]*kernel[2]+tmp[9661]*kernel[3]+tmp[9662]*kernel[4]+tmp[9663]*kernel[5]+tmp[9761]*kernel[6]+tmp[9762]*kernel[7]+tmp[9763]*kernel[8];
				ans[9663]<=tmp[9562]*kernel[0]+tmp[9563]*kernel[1]+tmp[9564]*kernel[2]+tmp[9662]*kernel[3]+tmp[9663]*kernel[4]+tmp[9664]*kernel[5]+tmp[9762]*kernel[6]+tmp[9763]*kernel[7]+tmp[9764]*kernel[8];
				ans[9664]<=tmp[9563]*kernel[0]+tmp[9564]*kernel[1]+tmp[9565]*kernel[2]+tmp[9663]*kernel[3]+tmp[9664]*kernel[4]+tmp[9665]*kernel[5]+tmp[9763]*kernel[6]+tmp[9764]*kernel[7]+tmp[9765]*kernel[8];
				ans[9665]<=tmp[9564]*kernel[0]+tmp[9565]*kernel[1]+tmp[9566]*kernel[2]+tmp[9664]*kernel[3]+tmp[9665]*kernel[4]+tmp[9666]*kernel[5]+tmp[9764]*kernel[6]+tmp[9765]*kernel[7]+tmp[9766]*kernel[8];
				ans[9666]<=tmp[9565]*kernel[0]+tmp[9566]*kernel[1]+tmp[9567]*kernel[2]+tmp[9665]*kernel[3]+tmp[9666]*kernel[4]+tmp[9667]*kernel[5]+tmp[9765]*kernel[6]+tmp[9766]*kernel[7]+tmp[9767]*kernel[8];
				ans[9667]<=tmp[9566]*kernel[0]+tmp[9567]*kernel[1]+tmp[9568]*kernel[2]+tmp[9666]*kernel[3]+tmp[9667]*kernel[4]+tmp[9668]*kernel[5]+tmp[9766]*kernel[6]+tmp[9767]*kernel[7]+tmp[9768]*kernel[8];
				ans[9668]<=tmp[9567]*kernel[0]+tmp[9568]*kernel[1]+tmp[9569]*kernel[2]+tmp[9667]*kernel[3]+tmp[9668]*kernel[4]+tmp[9669]*kernel[5]+tmp[9767]*kernel[6]+tmp[9768]*kernel[7]+tmp[9769]*kernel[8];
				ans[9669]<=tmp[9568]*kernel[0]+tmp[9569]*kernel[1]+tmp[9570]*kernel[2]+tmp[9668]*kernel[3]+tmp[9669]*kernel[4]+tmp[9670]*kernel[5]+tmp[9768]*kernel[6]+tmp[9769]*kernel[7]+tmp[9770]*kernel[8];
				ans[9670]<=tmp[9569]*kernel[0]+tmp[9570]*kernel[1]+tmp[9571]*kernel[2]+tmp[9669]*kernel[3]+tmp[9670]*kernel[4]+tmp[9671]*kernel[5]+tmp[9769]*kernel[6]+tmp[9770]*kernel[7]+tmp[9771]*kernel[8];
				ans[9671]<=tmp[9570]*kernel[0]+tmp[9571]*kernel[1]+tmp[9572]*kernel[2]+tmp[9670]*kernel[3]+tmp[9671]*kernel[4]+tmp[9672]*kernel[5]+tmp[9770]*kernel[6]+tmp[9771]*kernel[7]+tmp[9772]*kernel[8];
				ans[9672]<=tmp[9571]*kernel[0]+tmp[9572]*kernel[1]+tmp[9573]*kernel[2]+tmp[9671]*kernel[3]+tmp[9672]*kernel[4]+tmp[9673]*kernel[5]+tmp[9771]*kernel[6]+tmp[9772]*kernel[7]+tmp[9773]*kernel[8];
				ans[9673]<=tmp[9572]*kernel[0]+tmp[9573]*kernel[1]+tmp[9574]*kernel[2]+tmp[9672]*kernel[3]+tmp[9673]*kernel[4]+tmp[9674]*kernel[5]+tmp[9772]*kernel[6]+tmp[9773]*kernel[7]+tmp[9774]*kernel[8];
				ans[9674]<=tmp[9573]*kernel[0]+tmp[9574]*kernel[1]+tmp[9575]*kernel[2]+tmp[9673]*kernel[3]+tmp[9674]*kernel[4]+tmp[9675]*kernel[5]+tmp[9773]*kernel[6]+tmp[9774]*kernel[7]+tmp[9775]*kernel[8];
				ans[9675]<=tmp[9574]*kernel[0]+tmp[9575]*kernel[1]+tmp[9576]*kernel[2]+tmp[9674]*kernel[3]+tmp[9675]*kernel[4]+tmp[9676]*kernel[5]+tmp[9774]*kernel[6]+tmp[9775]*kernel[7]+tmp[9776]*kernel[8];
				ans[9676]<=tmp[9575]*kernel[0]+tmp[9576]*kernel[1]+tmp[9577]*kernel[2]+tmp[9675]*kernel[3]+tmp[9676]*kernel[4]+tmp[9677]*kernel[5]+tmp[9775]*kernel[6]+tmp[9776]*kernel[7]+tmp[9777]*kernel[8];
				ans[9677]<=tmp[9576]*kernel[0]+tmp[9577]*kernel[1]+tmp[9578]*kernel[2]+tmp[9676]*kernel[3]+tmp[9677]*kernel[4]+tmp[9678]*kernel[5]+tmp[9776]*kernel[6]+tmp[9777]*kernel[7]+tmp[9778]*kernel[8];
				ans[9678]<=tmp[9577]*kernel[0]+tmp[9578]*kernel[1]+tmp[9579]*kernel[2]+tmp[9677]*kernel[3]+tmp[9678]*kernel[4]+tmp[9679]*kernel[5]+tmp[9777]*kernel[6]+tmp[9778]*kernel[7]+tmp[9779]*kernel[8];
				ans[9679]<=tmp[9578]*kernel[0]+tmp[9579]*kernel[1]+tmp[9580]*kernel[2]+tmp[9678]*kernel[3]+tmp[9679]*kernel[4]+tmp[9680]*kernel[5]+tmp[9778]*kernel[6]+tmp[9779]*kernel[7]+tmp[9780]*kernel[8];
				ans[9680]<=tmp[9579]*kernel[0]+tmp[9580]*kernel[1]+tmp[9581]*kernel[2]+tmp[9679]*kernel[3]+tmp[9680]*kernel[4]+tmp[9681]*kernel[5]+tmp[9779]*kernel[6]+tmp[9780]*kernel[7]+tmp[9781]*kernel[8];
				ans[9681]<=tmp[9580]*kernel[0]+tmp[9581]*kernel[1]+tmp[9582]*kernel[2]+tmp[9680]*kernel[3]+tmp[9681]*kernel[4]+tmp[9682]*kernel[5]+tmp[9780]*kernel[6]+tmp[9781]*kernel[7]+tmp[9782]*kernel[8];
				ans[9682]<=tmp[9581]*kernel[0]+tmp[9582]*kernel[1]+tmp[9583]*kernel[2]+tmp[9681]*kernel[3]+tmp[9682]*kernel[4]+tmp[9683]*kernel[5]+tmp[9781]*kernel[6]+tmp[9782]*kernel[7]+tmp[9783]*kernel[8];
				ans[9683]<=tmp[9582]*kernel[0]+tmp[9583]*kernel[1]+tmp[9584]*kernel[2]+tmp[9682]*kernel[3]+tmp[9683]*kernel[4]+tmp[9684]*kernel[5]+tmp[9782]*kernel[6]+tmp[9783]*kernel[7]+tmp[9784]*kernel[8];
				ans[9684]<=tmp[9583]*kernel[0]+tmp[9584]*kernel[1]+tmp[9585]*kernel[2]+tmp[9683]*kernel[3]+tmp[9684]*kernel[4]+tmp[9685]*kernel[5]+tmp[9783]*kernel[6]+tmp[9784]*kernel[7]+tmp[9785]*kernel[8];
				ans[9685]<=tmp[9584]*kernel[0]+tmp[9585]*kernel[1]+tmp[9586]*kernel[2]+tmp[9684]*kernel[3]+tmp[9685]*kernel[4]+tmp[9686]*kernel[5]+tmp[9784]*kernel[6]+tmp[9785]*kernel[7]+tmp[9786]*kernel[8];
				ans[9686]<=tmp[9585]*kernel[0]+tmp[9586]*kernel[1]+tmp[9587]*kernel[2]+tmp[9685]*kernel[3]+tmp[9686]*kernel[4]+tmp[9687]*kernel[5]+tmp[9785]*kernel[6]+tmp[9786]*kernel[7]+tmp[9787]*kernel[8];
				ans[9687]<=tmp[9586]*kernel[0]+tmp[9587]*kernel[1]+tmp[9588]*kernel[2]+tmp[9686]*kernel[3]+tmp[9687]*kernel[4]+tmp[9688]*kernel[5]+tmp[9786]*kernel[6]+tmp[9787]*kernel[7]+tmp[9788]*kernel[8];
				ans[9688]<=tmp[9587]*kernel[0]+tmp[9588]*kernel[1]+tmp[9589]*kernel[2]+tmp[9687]*kernel[3]+tmp[9688]*kernel[4]+tmp[9689]*kernel[5]+tmp[9787]*kernel[6]+tmp[9788]*kernel[7]+tmp[9789]*kernel[8];
				ans[9689]<=tmp[9588]*kernel[0]+tmp[9589]*kernel[1]+tmp[9590]*kernel[2]+tmp[9688]*kernel[3]+tmp[9689]*kernel[4]+tmp[9690]*kernel[5]+tmp[9788]*kernel[6]+tmp[9789]*kernel[7]+tmp[9790]*kernel[8];
				ans[9690]<=tmp[9589]*kernel[0]+tmp[9590]*kernel[1]+tmp[9591]*kernel[2]+tmp[9689]*kernel[3]+tmp[9690]*kernel[4]+tmp[9691]*kernel[5]+tmp[9789]*kernel[6]+tmp[9790]*kernel[7]+tmp[9791]*kernel[8];
				ans[9691]<=tmp[9590]*kernel[0]+tmp[9591]*kernel[1]+tmp[9592]*kernel[2]+tmp[9690]*kernel[3]+tmp[9691]*kernel[4]+tmp[9692]*kernel[5]+tmp[9790]*kernel[6]+tmp[9791]*kernel[7]+tmp[9792]*kernel[8];
				ans[9692]<=tmp[9591]*kernel[0]+tmp[9592]*kernel[1]+tmp[9593]*kernel[2]+tmp[9691]*kernel[3]+tmp[9692]*kernel[4]+tmp[9693]*kernel[5]+tmp[9791]*kernel[6]+tmp[9792]*kernel[7]+tmp[9793]*kernel[8];
				ans[9693]<=tmp[9592]*kernel[0]+tmp[9593]*kernel[1]+tmp[9594]*kernel[2]+tmp[9692]*kernel[3]+tmp[9693]*kernel[4]+tmp[9694]*kernel[5]+tmp[9792]*kernel[6]+tmp[9793]*kernel[7]+tmp[9794]*kernel[8];
				ans[9694]<=tmp[9593]*kernel[0]+tmp[9594]*kernel[1]+tmp[9595]*kernel[2]+tmp[9693]*kernel[3]+tmp[9694]*kernel[4]+tmp[9695]*kernel[5]+tmp[9793]*kernel[6]+tmp[9794]*kernel[7]+tmp[9795]*kernel[8];
				ans[9695]<=tmp[9594]*kernel[0]+tmp[9595]*kernel[1]+tmp[9596]*kernel[2]+tmp[9694]*kernel[3]+tmp[9695]*kernel[4]+tmp[9696]*kernel[5]+tmp[9794]*kernel[6]+tmp[9795]*kernel[7]+tmp[9796]*kernel[8];
				ans[9696]<=tmp[9595]*kernel[0]+tmp[9596]*kernel[1]+tmp[9597]*kernel[2]+tmp[9695]*kernel[3]+tmp[9696]*kernel[4]+tmp[9697]*kernel[5]+tmp[9795]*kernel[6]+tmp[9796]*kernel[7]+tmp[9797]*kernel[8];
				ans[9697]<=tmp[9596]*kernel[0]+tmp[9597]*kernel[1]+tmp[9598]*kernel[2]+tmp[9696]*kernel[3]+tmp[9697]*kernel[4]+tmp[9698]*kernel[5]+tmp[9796]*kernel[6]+tmp[9797]*kernel[7]+tmp[9798]*kernel[8];
				ans[9698]<=tmp[9597]*kernel[0]+tmp[9598]*kernel[1]+tmp[9599]*kernel[2]+tmp[9697]*kernel[3]+tmp[9698]*kernel[4]+tmp[9699]*kernel[5]+tmp[9797]*kernel[6]+tmp[9798]*kernel[7]+tmp[9799]*kernel[8];
				ans[9699]<=tmp[9598]*kernel[0]+tmp[9599]*kernel[1]+tmp[9698]*kernel[3]+tmp[9699]*kernel[4]+tmp[9798]*kernel[6]+tmp[9799]*kernel[7];
				ans[9700]<=tmp[9600]*kernel[1]+tmp[9601]*kernel[2]+tmp[9700]*kernel[4]+tmp[9701]*kernel[5]+tmp[9800]*kernel[7]+tmp[9801]*kernel[8];
				ans[9701]<=tmp[9600]*kernel[0]+tmp[9601]*kernel[1]+tmp[9602]*kernel[2]+tmp[9700]*kernel[3]+tmp[9701]*kernel[4]+tmp[9702]*kernel[5]+tmp[9800]*kernel[6]+tmp[9801]*kernel[7]+tmp[9802]*kernel[8];
				ans[9702]<=tmp[9601]*kernel[0]+tmp[9602]*kernel[1]+tmp[9603]*kernel[2]+tmp[9701]*kernel[3]+tmp[9702]*kernel[4]+tmp[9703]*kernel[5]+tmp[9801]*kernel[6]+tmp[9802]*kernel[7]+tmp[9803]*kernel[8];
				ans[9703]<=tmp[9602]*kernel[0]+tmp[9603]*kernel[1]+tmp[9604]*kernel[2]+tmp[9702]*kernel[3]+tmp[9703]*kernel[4]+tmp[9704]*kernel[5]+tmp[9802]*kernel[6]+tmp[9803]*kernel[7]+tmp[9804]*kernel[8];
				ans[9704]<=tmp[9603]*kernel[0]+tmp[9604]*kernel[1]+tmp[9605]*kernel[2]+tmp[9703]*kernel[3]+tmp[9704]*kernel[4]+tmp[9705]*kernel[5]+tmp[9803]*kernel[6]+tmp[9804]*kernel[7]+tmp[9805]*kernel[8];
				ans[9705]<=tmp[9604]*kernel[0]+tmp[9605]*kernel[1]+tmp[9606]*kernel[2]+tmp[9704]*kernel[3]+tmp[9705]*kernel[4]+tmp[9706]*kernel[5]+tmp[9804]*kernel[6]+tmp[9805]*kernel[7]+tmp[9806]*kernel[8];
				ans[9706]<=tmp[9605]*kernel[0]+tmp[9606]*kernel[1]+tmp[9607]*kernel[2]+tmp[9705]*kernel[3]+tmp[9706]*kernel[4]+tmp[9707]*kernel[5]+tmp[9805]*kernel[6]+tmp[9806]*kernel[7]+tmp[9807]*kernel[8];
				ans[9707]<=tmp[9606]*kernel[0]+tmp[9607]*kernel[1]+tmp[9608]*kernel[2]+tmp[9706]*kernel[3]+tmp[9707]*kernel[4]+tmp[9708]*kernel[5]+tmp[9806]*kernel[6]+tmp[9807]*kernel[7]+tmp[9808]*kernel[8];
				ans[9708]<=tmp[9607]*kernel[0]+tmp[9608]*kernel[1]+tmp[9609]*kernel[2]+tmp[9707]*kernel[3]+tmp[9708]*kernel[4]+tmp[9709]*kernel[5]+tmp[9807]*kernel[6]+tmp[9808]*kernel[7]+tmp[9809]*kernel[8];
				ans[9709]<=tmp[9608]*kernel[0]+tmp[9609]*kernel[1]+tmp[9610]*kernel[2]+tmp[9708]*kernel[3]+tmp[9709]*kernel[4]+tmp[9710]*kernel[5]+tmp[9808]*kernel[6]+tmp[9809]*kernel[7]+tmp[9810]*kernel[8];
				ans[9710]<=tmp[9609]*kernel[0]+tmp[9610]*kernel[1]+tmp[9611]*kernel[2]+tmp[9709]*kernel[3]+tmp[9710]*kernel[4]+tmp[9711]*kernel[5]+tmp[9809]*kernel[6]+tmp[9810]*kernel[7]+tmp[9811]*kernel[8];
				ans[9711]<=tmp[9610]*kernel[0]+tmp[9611]*kernel[1]+tmp[9612]*kernel[2]+tmp[9710]*kernel[3]+tmp[9711]*kernel[4]+tmp[9712]*kernel[5]+tmp[9810]*kernel[6]+tmp[9811]*kernel[7]+tmp[9812]*kernel[8];
				ans[9712]<=tmp[9611]*kernel[0]+tmp[9612]*kernel[1]+tmp[9613]*kernel[2]+tmp[9711]*kernel[3]+tmp[9712]*kernel[4]+tmp[9713]*kernel[5]+tmp[9811]*kernel[6]+tmp[9812]*kernel[7]+tmp[9813]*kernel[8];
				ans[9713]<=tmp[9612]*kernel[0]+tmp[9613]*kernel[1]+tmp[9614]*kernel[2]+tmp[9712]*kernel[3]+tmp[9713]*kernel[4]+tmp[9714]*kernel[5]+tmp[9812]*kernel[6]+tmp[9813]*kernel[7]+tmp[9814]*kernel[8];
				ans[9714]<=tmp[9613]*kernel[0]+tmp[9614]*kernel[1]+tmp[9615]*kernel[2]+tmp[9713]*kernel[3]+tmp[9714]*kernel[4]+tmp[9715]*kernel[5]+tmp[9813]*kernel[6]+tmp[9814]*kernel[7]+tmp[9815]*kernel[8];
				ans[9715]<=tmp[9614]*kernel[0]+tmp[9615]*kernel[1]+tmp[9616]*kernel[2]+tmp[9714]*kernel[3]+tmp[9715]*kernel[4]+tmp[9716]*kernel[5]+tmp[9814]*kernel[6]+tmp[9815]*kernel[7]+tmp[9816]*kernel[8];
				ans[9716]<=tmp[9615]*kernel[0]+tmp[9616]*kernel[1]+tmp[9617]*kernel[2]+tmp[9715]*kernel[3]+tmp[9716]*kernel[4]+tmp[9717]*kernel[5]+tmp[9815]*kernel[6]+tmp[9816]*kernel[7]+tmp[9817]*kernel[8];
				ans[9717]<=tmp[9616]*kernel[0]+tmp[9617]*kernel[1]+tmp[9618]*kernel[2]+tmp[9716]*kernel[3]+tmp[9717]*kernel[4]+tmp[9718]*kernel[5]+tmp[9816]*kernel[6]+tmp[9817]*kernel[7]+tmp[9818]*kernel[8];
				ans[9718]<=tmp[9617]*kernel[0]+tmp[9618]*kernel[1]+tmp[9619]*kernel[2]+tmp[9717]*kernel[3]+tmp[9718]*kernel[4]+tmp[9719]*kernel[5]+tmp[9817]*kernel[6]+tmp[9818]*kernel[7]+tmp[9819]*kernel[8];
				ans[9719]<=tmp[9618]*kernel[0]+tmp[9619]*kernel[1]+tmp[9620]*kernel[2]+tmp[9718]*kernel[3]+tmp[9719]*kernel[4]+tmp[9720]*kernel[5]+tmp[9818]*kernel[6]+tmp[9819]*kernel[7]+tmp[9820]*kernel[8];
				ans[9720]<=tmp[9619]*kernel[0]+tmp[9620]*kernel[1]+tmp[9621]*kernel[2]+tmp[9719]*kernel[3]+tmp[9720]*kernel[4]+tmp[9721]*kernel[5]+tmp[9819]*kernel[6]+tmp[9820]*kernel[7]+tmp[9821]*kernel[8];
				ans[9721]<=tmp[9620]*kernel[0]+tmp[9621]*kernel[1]+tmp[9622]*kernel[2]+tmp[9720]*kernel[3]+tmp[9721]*kernel[4]+tmp[9722]*kernel[5]+tmp[9820]*kernel[6]+tmp[9821]*kernel[7]+tmp[9822]*kernel[8];
				ans[9722]<=tmp[9621]*kernel[0]+tmp[9622]*kernel[1]+tmp[9623]*kernel[2]+tmp[9721]*kernel[3]+tmp[9722]*kernel[4]+tmp[9723]*kernel[5]+tmp[9821]*kernel[6]+tmp[9822]*kernel[7]+tmp[9823]*kernel[8];
				ans[9723]<=tmp[9622]*kernel[0]+tmp[9623]*kernel[1]+tmp[9624]*kernel[2]+tmp[9722]*kernel[3]+tmp[9723]*kernel[4]+tmp[9724]*kernel[5]+tmp[9822]*kernel[6]+tmp[9823]*kernel[7]+tmp[9824]*kernel[8];
				ans[9724]<=tmp[9623]*kernel[0]+tmp[9624]*kernel[1]+tmp[9625]*kernel[2]+tmp[9723]*kernel[3]+tmp[9724]*kernel[4]+tmp[9725]*kernel[5]+tmp[9823]*kernel[6]+tmp[9824]*kernel[7]+tmp[9825]*kernel[8];
				ans[9725]<=tmp[9624]*kernel[0]+tmp[9625]*kernel[1]+tmp[9626]*kernel[2]+tmp[9724]*kernel[3]+tmp[9725]*kernel[4]+tmp[9726]*kernel[5]+tmp[9824]*kernel[6]+tmp[9825]*kernel[7]+tmp[9826]*kernel[8];
				ans[9726]<=tmp[9625]*kernel[0]+tmp[9626]*kernel[1]+tmp[9627]*kernel[2]+tmp[9725]*kernel[3]+tmp[9726]*kernel[4]+tmp[9727]*kernel[5]+tmp[9825]*kernel[6]+tmp[9826]*kernel[7]+tmp[9827]*kernel[8];
				ans[9727]<=tmp[9626]*kernel[0]+tmp[9627]*kernel[1]+tmp[9628]*kernel[2]+tmp[9726]*kernel[3]+tmp[9727]*kernel[4]+tmp[9728]*kernel[5]+tmp[9826]*kernel[6]+tmp[9827]*kernel[7]+tmp[9828]*kernel[8];
				ans[9728]<=tmp[9627]*kernel[0]+tmp[9628]*kernel[1]+tmp[9629]*kernel[2]+tmp[9727]*kernel[3]+tmp[9728]*kernel[4]+tmp[9729]*kernel[5]+tmp[9827]*kernel[6]+tmp[9828]*kernel[7]+tmp[9829]*kernel[8];
				ans[9729]<=tmp[9628]*kernel[0]+tmp[9629]*kernel[1]+tmp[9630]*kernel[2]+tmp[9728]*kernel[3]+tmp[9729]*kernel[4]+tmp[9730]*kernel[5]+tmp[9828]*kernel[6]+tmp[9829]*kernel[7]+tmp[9830]*kernel[8];
				ans[9730]<=tmp[9629]*kernel[0]+tmp[9630]*kernel[1]+tmp[9631]*kernel[2]+tmp[9729]*kernel[3]+tmp[9730]*kernel[4]+tmp[9731]*kernel[5]+tmp[9829]*kernel[6]+tmp[9830]*kernel[7]+tmp[9831]*kernel[8];
				ans[9731]<=tmp[9630]*kernel[0]+tmp[9631]*kernel[1]+tmp[9632]*kernel[2]+tmp[9730]*kernel[3]+tmp[9731]*kernel[4]+tmp[9732]*kernel[5]+tmp[9830]*kernel[6]+tmp[9831]*kernel[7]+tmp[9832]*kernel[8];
				ans[9732]<=tmp[9631]*kernel[0]+tmp[9632]*kernel[1]+tmp[9633]*kernel[2]+tmp[9731]*kernel[3]+tmp[9732]*kernel[4]+tmp[9733]*kernel[5]+tmp[9831]*kernel[6]+tmp[9832]*kernel[7]+tmp[9833]*kernel[8];
				ans[9733]<=tmp[9632]*kernel[0]+tmp[9633]*kernel[1]+tmp[9634]*kernel[2]+tmp[9732]*kernel[3]+tmp[9733]*kernel[4]+tmp[9734]*kernel[5]+tmp[9832]*kernel[6]+tmp[9833]*kernel[7]+tmp[9834]*kernel[8];
				ans[9734]<=tmp[9633]*kernel[0]+tmp[9634]*kernel[1]+tmp[9635]*kernel[2]+tmp[9733]*kernel[3]+tmp[9734]*kernel[4]+tmp[9735]*kernel[5]+tmp[9833]*kernel[6]+tmp[9834]*kernel[7]+tmp[9835]*kernel[8];
				ans[9735]<=tmp[9634]*kernel[0]+tmp[9635]*kernel[1]+tmp[9636]*kernel[2]+tmp[9734]*kernel[3]+tmp[9735]*kernel[4]+tmp[9736]*kernel[5]+tmp[9834]*kernel[6]+tmp[9835]*kernel[7]+tmp[9836]*kernel[8];
				ans[9736]<=tmp[9635]*kernel[0]+tmp[9636]*kernel[1]+tmp[9637]*kernel[2]+tmp[9735]*kernel[3]+tmp[9736]*kernel[4]+tmp[9737]*kernel[5]+tmp[9835]*kernel[6]+tmp[9836]*kernel[7]+tmp[9837]*kernel[8];
				ans[9737]<=tmp[9636]*kernel[0]+tmp[9637]*kernel[1]+tmp[9638]*kernel[2]+tmp[9736]*kernel[3]+tmp[9737]*kernel[4]+tmp[9738]*kernel[5]+tmp[9836]*kernel[6]+tmp[9837]*kernel[7]+tmp[9838]*kernel[8];
				ans[9738]<=tmp[9637]*kernel[0]+tmp[9638]*kernel[1]+tmp[9639]*kernel[2]+tmp[9737]*kernel[3]+tmp[9738]*kernel[4]+tmp[9739]*kernel[5]+tmp[9837]*kernel[6]+tmp[9838]*kernel[7]+tmp[9839]*kernel[8];
				ans[9739]<=tmp[9638]*kernel[0]+tmp[9639]*kernel[1]+tmp[9640]*kernel[2]+tmp[9738]*kernel[3]+tmp[9739]*kernel[4]+tmp[9740]*kernel[5]+tmp[9838]*kernel[6]+tmp[9839]*kernel[7]+tmp[9840]*kernel[8];
				ans[9740]<=tmp[9639]*kernel[0]+tmp[9640]*kernel[1]+tmp[9641]*kernel[2]+tmp[9739]*kernel[3]+tmp[9740]*kernel[4]+tmp[9741]*kernel[5]+tmp[9839]*kernel[6]+tmp[9840]*kernel[7]+tmp[9841]*kernel[8];
				ans[9741]<=tmp[9640]*kernel[0]+tmp[9641]*kernel[1]+tmp[9642]*kernel[2]+tmp[9740]*kernel[3]+tmp[9741]*kernel[4]+tmp[9742]*kernel[5]+tmp[9840]*kernel[6]+tmp[9841]*kernel[7]+tmp[9842]*kernel[8];
				ans[9742]<=tmp[9641]*kernel[0]+tmp[9642]*kernel[1]+tmp[9643]*kernel[2]+tmp[9741]*kernel[3]+tmp[9742]*kernel[4]+tmp[9743]*kernel[5]+tmp[9841]*kernel[6]+tmp[9842]*kernel[7]+tmp[9843]*kernel[8];
				ans[9743]<=tmp[9642]*kernel[0]+tmp[9643]*kernel[1]+tmp[9644]*kernel[2]+tmp[9742]*kernel[3]+tmp[9743]*kernel[4]+tmp[9744]*kernel[5]+tmp[9842]*kernel[6]+tmp[9843]*kernel[7]+tmp[9844]*kernel[8];
				ans[9744]<=tmp[9643]*kernel[0]+tmp[9644]*kernel[1]+tmp[9645]*kernel[2]+tmp[9743]*kernel[3]+tmp[9744]*kernel[4]+tmp[9745]*kernel[5]+tmp[9843]*kernel[6]+tmp[9844]*kernel[7]+tmp[9845]*kernel[8];
				ans[9745]<=tmp[9644]*kernel[0]+tmp[9645]*kernel[1]+tmp[9646]*kernel[2]+tmp[9744]*kernel[3]+tmp[9745]*kernel[4]+tmp[9746]*kernel[5]+tmp[9844]*kernel[6]+tmp[9845]*kernel[7]+tmp[9846]*kernel[8];
				ans[9746]<=tmp[9645]*kernel[0]+tmp[9646]*kernel[1]+tmp[9647]*kernel[2]+tmp[9745]*kernel[3]+tmp[9746]*kernel[4]+tmp[9747]*kernel[5]+tmp[9845]*kernel[6]+tmp[9846]*kernel[7]+tmp[9847]*kernel[8];
				ans[9747]<=tmp[9646]*kernel[0]+tmp[9647]*kernel[1]+tmp[9648]*kernel[2]+tmp[9746]*kernel[3]+tmp[9747]*kernel[4]+tmp[9748]*kernel[5]+tmp[9846]*kernel[6]+tmp[9847]*kernel[7]+tmp[9848]*kernel[8];
				ans[9748]<=tmp[9647]*kernel[0]+tmp[9648]*kernel[1]+tmp[9649]*kernel[2]+tmp[9747]*kernel[3]+tmp[9748]*kernel[4]+tmp[9749]*kernel[5]+tmp[9847]*kernel[6]+tmp[9848]*kernel[7]+tmp[9849]*kernel[8];
				ans[9749]<=tmp[9648]*kernel[0]+tmp[9649]*kernel[1]+tmp[9650]*kernel[2]+tmp[9748]*kernel[3]+tmp[9749]*kernel[4]+tmp[9750]*kernel[5]+tmp[9848]*kernel[6]+tmp[9849]*kernel[7]+tmp[9850]*kernel[8];
				ans[9750]<=tmp[9649]*kernel[0]+tmp[9650]*kernel[1]+tmp[9651]*kernel[2]+tmp[9749]*kernel[3]+tmp[9750]*kernel[4]+tmp[9751]*kernel[5]+tmp[9849]*kernel[6]+tmp[9850]*kernel[7]+tmp[9851]*kernel[8];
				ans[9751]<=tmp[9650]*kernel[0]+tmp[9651]*kernel[1]+tmp[9652]*kernel[2]+tmp[9750]*kernel[3]+tmp[9751]*kernel[4]+tmp[9752]*kernel[5]+tmp[9850]*kernel[6]+tmp[9851]*kernel[7]+tmp[9852]*kernel[8];
				ans[9752]<=tmp[9651]*kernel[0]+tmp[9652]*kernel[1]+tmp[9653]*kernel[2]+tmp[9751]*kernel[3]+tmp[9752]*kernel[4]+tmp[9753]*kernel[5]+tmp[9851]*kernel[6]+tmp[9852]*kernel[7]+tmp[9853]*kernel[8];
				ans[9753]<=tmp[9652]*kernel[0]+tmp[9653]*kernel[1]+tmp[9654]*kernel[2]+tmp[9752]*kernel[3]+tmp[9753]*kernel[4]+tmp[9754]*kernel[5]+tmp[9852]*kernel[6]+tmp[9853]*kernel[7]+tmp[9854]*kernel[8];
				ans[9754]<=tmp[9653]*kernel[0]+tmp[9654]*kernel[1]+tmp[9655]*kernel[2]+tmp[9753]*kernel[3]+tmp[9754]*kernel[4]+tmp[9755]*kernel[5]+tmp[9853]*kernel[6]+tmp[9854]*kernel[7]+tmp[9855]*kernel[8];
				ans[9755]<=tmp[9654]*kernel[0]+tmp[9655]*kernel[1]+tmp[9656]*kernel[2]+tmp[9754]*kernel[3]+tmp[9755]*kernel[4]+tmp[9756]*kernel[5]+tmp[9854]*kernel[6]+tmp[9855]*kernel[7]+tmp[9856]*kernel[8];
				ans[9756]<=tmp[9655]*kernel[0]+tmp[9656]*kernel[1]+tmp[9657]*kernel[2]+tmp[9755]*kernel[3]+tmp[9756]*kernel[4]+tmp[9757]*kernel[5]+tmp[9855]*kernel[6]+tmp[9856]*kernel[7]+tmp[9857]*kernel[8];
				ans[9757]<=tmp[9656]*kernel[0]+tmp[9657]*kernel[1]+tmp[9658]*kernel[2]+tmp[9756]*kernel[3]+tmp[9757]*kernel[4]+tmp[9758]*kernel[5]+tmp[9856]*kernel[6]+tmp[9857]*kernel[7]+tmp[9858]*kernel[8];
				ans[9758]<=tmp[9657]*kernel[0]+tmp[9658]*kernel[1]+tmp[9659]*kernel[2]+tmp[9757]*kernel[3]+tmp[9758]*kernel[4]+tmp[9759]*kernel[5]+tmp[9857]*kernel[6]+tmp[9858]*kernel[7]+tmp[9859]*kernel[8];
				ans[9759]<=tmp[9658]*kernel[0]+tmp[9659]*kernel[1]+tmp[9660]*kernel[2]+tmp[9758]*kernel[3]+tmp[9759]*kernel[4]+tmp[9760]*kernel[5]+tmp[9858]*kernel[6]+tmp[9859]*kernel[7]+tmp[9860]*kernel[8];
				ans[9760]<=tmp[9659]*kernel[0]+tmp[9660]*kernel[1]+tmp[9661]*kernel[2]+tmp[9759]*kernel[3]+tmp[9760]*kernel[4]+tmp[9761]*kernel[5]+tmp[9859]*kernel[6]+tmp[9860]*kernel[7]+tmp[9861]*kernel[8];
				ans[9761]<=tmp[9660]*kernel[0]+tmp[9661]*kernel[1]+tmp[9662]*kernel[2]+tmp[9760]*kernel[3]+tmp[9761]*kernel[4]+tmp[9762]*kernel[5]+tmp[9860]*kernel[6]+tmp[9861]*kernel[7]+tmp[9862]*kernel[8];
				ans[9762]<=tmp[9661]*kernel[0]+tmp[9662]*kernel[1]+tmp[9663]*kernel[2]+tmp[9761]*kernel[3]+tmp[9762]*kernel[4]+tmp[9763]*kernel[5]+tmp[9861]*kernel[6]+tmp[9862]*kernel[7]+tmp[9863]*kernel[8];
				ans[9763]<=tmp[9662]*kernel[0]+tmp[9663]*kernel[1]+tmp[9664]*kernel[2]+tmp[9762]*kernel[3]+tmp[9763]*kernel[4]+tmp[9764]*kernel[5]+tmp[9862]*kernel[6]+tmp[9863]*kernel[7]+tmp[9864]*kernel[8];
				ans[9764]<=tmp[9663]*kernel[0]+tmp[9664]*kernel[1]+tmp[9665]*kernel[2]+tmp[9763]*kernel[3]+tmp[9764]*kernel[4]+tmp[9765]*kernel[5]+tmp[9863]*kernel[6]+tmp[9864]*kernel[7]+tmp[9865]*kernel[8];
				ans[9765]<=tmp[9664]*kernel[0]+tmp[9665]*kernel[1]+tmp[9666]*kernel[2]+tmp[9764]*kernel[3]+tmp[9765]*kernel[4]+tmp[9766]*kernel[5]+tmp[9864]*kernel[6]+tmp[9865]*kernel[7]+tmp[9866]*kernel[8];
				ans[9766]<=tmp[9665]*kernel[0]+tmp[9666]*kernel[1]+tmp[9667]*kernel[2]+tmp[9765]*kernel[3]+tmp[9766]*kernel[4]+tmp[9767]*kernel[5]+tmp[9865]*kernel[6]+tmp[9866]*kernel[7]+tmp[9867]*kernel[8];
				ans[9767]<=tmp[9666]*kernel[0]+tmp[9667]*kernel[1]+tmp[9668]*kernel[2]+tmp[9766]*kernel[3]+tmp[9767]*kernel[4]+tmp[9768]*kernel[5]+tmp[9866]*kernel[6]+tmp[9867]*kernel[7]+tmp[9868]*kernel[8];
				ans[9768]<=tmp[9667]*kernel[0]+tmp[9668]*kernel[1]+tmp[9669]*kernel[2]+tmp[9767]*kernel[3]+tmp[9768]*kernel[4]+tmp[9769]*kernel[5]+tmp[9867]*kernel[6]+tmp[9868]*kernel[7]+tmp[9869]*kernel[8];
				ans[9769]<=tmp[9668]*kernel[0]+tmp[9669]*kernel[1]+tmp[9670]*kernel[2]+tmp[9768]*kernel[3]+tmp[9769]*kernel[4]+tmp[9770]*kernel[5]+tmp[9868]*kernel[6]+tmp[9869]*kernel[7]+tmp[9870]*kernel[8];
				ans[9770]<=tmp[9669]*kernel[0]+tmp[9670]*kernel[1]+tmp[9671]*kernel[2]+tmp[9769]*kernel[3]+tmp[9770]*kernel[4]+tmp[9771]*kernel[5]+tmp[9869]*kernel[6]+tmp[9870]*kernel[7]+tmp[9871]*kernel[8];
				ans[9771]<=tmp[9670]*kernel[0]+tmp[9671]*kernel[1]+tmp[9672]*kernel[2]+tmp[9770]*kernel[3]+tmp[9771]*kernel[4]+tmp[9772]*kernel[5]+tmp[9870]*kernel[6]+tmp[9871]*kernel[7]+tmp[9872]*kernel[8];
				ans[9772]<=tmp[9671]*kernel[0]+tmp[9672]*kernel[1]+tmp[9673]*kernel[2]+tmp[9771]*kernel[3]+tmp[9772]*kernel[4]+tmp[9773]*kernel[5]+tmp[9871]*kernel[6]+tmp[9872]*kernel[7]+tmp[9873]*kernel[8];
				ans[9773]<=tmp[9672]*kernel[0]+tmp[9673]*kernel[1]+tmp[9674]*kernel[2]+tmp[9772]*kernel[3]+tmp[9773]*kernel[4]+tmp[9774]*kernel[5]+tmp[9872]*kernel[6]+tmp[9873]*kernel[7]+tmp[9874]*kernel[8];
				ans[9774]<=tmp[9673]*kernel[0]+tmp[9674]*kernel[1]+tmp[9675]*kernel[2]+tmp[9773]*kernel[3]+tmp[9774]*kernel[4]+tmp[9775]*kernel[5]+tmp[9873]*kernel[6]+tmp[9874]*kernel[7]+tmp[9875]*kernel[8];
				ans[9775]<=tmp[9674]*kernel[0]+tmp[9675]*kernel[1]+tmp[9676]*kernel[2]+tmp[9774]*kernel[3]+tmp[9775]*kernel[4]+tmp[9776]*kernel[5]+tmp[9874]*kernel[6]+tmp[9875]*kernel[7]+tmp[9876]*kernel[8];
				ans[9776]<=tmp[9675]*kernel[0]+tmp[9676]*kernel[1]+tmp[9677]*kernel[2]+tmp[9775]*kernel[3]+tmp[9776]*kernel[4]+tmp[9777]*kernel[5]+tmp[9875]*kernel[6]+tmp[9876]*kernel[7]+tmp[9877]*kernel[8];
				ans[9777]<=tmp[9676]*kernel[0]+tmp[9677]*kernel[1]+tmp[9678]*kernel[2]+tmp[9776]*kernel[3]+tmp[9777]*kernel[4]+tmp[9778]*kernel[5]+tmp[9876]*kernel[6]+tmp[9877]*kernel[7]+tmp[9878]*kernel[8];
				ans[9778]<=tmp[9677]*kernel[0]+tmp[9678]*kernel[1]+tmp[9679]*kernel[2]+tmp[9777]*kernel[3]+tmp[9778]*kernel[4]+tmp[9779]*kernel[5]+tmp[9877]*kernel[6]+tmp[9878]*kernel[7]+tmp[9879]*kernel[8];
				ans[9779]<=tmp[9678]*kernel[0]+tmp[9679]*kernel[1]+tmp[9680]*kernel[2]+tmp[9778]*kernel[3]+tmp[9779]*kernel[4]+tmp[9780]*kernel[5]+tmp[9878]*kernel[6]+tmp[9879]*kernel[7]+tmp[9880]*kernel[8];
				ans[9780]<=tmp[9679]*kernel[0]+tmp[9680]*kernel[1]+tmp[9681]*kernel[2]+tmp[9779]*kernel[3]+tmp[9780]*kernel[4]+tmp[9781]*kernel[5]+tmp[9879]*kernel[6]+tmp[9880]*kernel[7]+tmp[9881]*kernel[8];
				ans[9781]<=tmp[9680]*kernel[0]+tmp[9681]*kernel[1]+tmp[9682]*kernel[2]+tmp[9780]*kernel[3]+tmp[9781]*kernel[4]+tmp[9782]*kernel[5]+tmp[9880]*kernel[6]+tmp[9881]*kernel[7]+tmp[9882]*kernel[8];
				ans[9782]<=tmp[9681]*kernel[0]+tmp[9682]*kernel[1]+tmp[9683]*kernel[2]+tmp[9781]*kernel[3]+tmp[9782]*kernel[4]+tmp[9783]*kernel[5]+tmp[9881]*kernel[6]+tmp[9882]*kernel[7]+tmp[9883]*kernel[8];
				ans[9783]<=tmp[9682]*kernel[0]+tmp[9683]*kernel[1]+tmp[9684]*kernel[2]+tmp[9782]*kernel[3]+tmp[9783]*kernel[4]+tmp[9784]*kernel[5]+tmp[9882]*kernel[6]+tmp[9883]*kernel[7]+tmp[9884]*kernel[8];
				ans[9784]<=tmp[9683]*kernel[0]+tmp[9684]*kernel[1]+tmp[9685]*kernel[2]+tmp[9783]*kernel[3]+tmp[9784]*kernel[4]+tmp[9785]*kernel[5]+tmp[9883]*kernel[6]+tmp[9884]*kernel[7]+tmp[9885]*kernel[8];
				ans[9785]<=tmp[9684]*kernel[0]+tmp[9685]*kernel[1]+tmp[9686]*kernel[2]+tmp[9784]*kernel[3]+tmp[9785]*kernel[4]+tmp[9786]*kernel[5]+tmp[9884]*kernel[6]+tmp[9885]*kernel[7]+tmp[9886]*kernel[8];
				ans[9786]<=tmp[9685]*kernel[0]+tmp[9686]*kernel[1]+tmp[9687]*kernel[2]+tmp[9785]*kernel[3]+tmp[9786]*kernel[4]+tmp[9787]*kernel[5]+tmp[9885]*kernel[6]+tmp[9886]*kernel[7]+tmp[9887]*kernel[8];
				ans[9787]<=tmp[9686]*kernel[0]+tmp[9687]*kernel[1]+tmp[9688]*kernel[2]+tmp[9786]*kernel[3]+tmp[9787]*kernel[4]+tmp[9788]*kernel[5]+tmp[9886]*kernel[6]+tmp[9887]*kernel[7]+tmp[9888]*kernel[8];
				ans[9788]<=tmp[9687]*kernel[0]+tmp[9688]*kernel[1]+tmp[9689]*kernel[2]+tmp[9787]*kernel[3]+tmp[9788]*kernel[4]+tmp[9789]*kernel[5]+tmp[9887]*kernel[6]+tmp[9888]*kernel[7]+tmp[9889]*kernel[8];
				ans[9789]<=tmp[9688]*kernel[0]+tmp[9689]*kernel[1]+tmp[9690]*kernel[2]+tmp[9788]*kernel[3]+tmp[9789]*kernel[4]+tmp[9790]*kernel[5]+tmp[9888]*kernel[6]+tmp[9889]*kernel[7]+tmp[9890]*kernel[8];
				ans[9790]<=tmp[9689]*kernel[0]+tmp[9690]*kernel[1]+tmp[9691]*kernel[2]+tmp[9789]*kernel[3]+tmp[9790]*kernel[4]+tmp[9791]*kernel[5]+tmp[9889]*kernel[6]+tmp[9890]*kernel[7]+tmp[9891]*kernel[8];
				ans[9791]<=tmp[9690]*kernel[0]+tmp[9691]*kernel[1]+tmp[9692]*kernel[2]+tmp[9790]*kernel[3]+tmp[9791]*kernel[4]+tmp[9792]*kernel[5]+tmp[9890]*kernel[6]+tmp[9891]*kernel[7]+tmp[9892]*kernel[8];
				ans[9792]<=tmp[9691]*kernel[0]+tmp[9692]*kernel[1]+tmp[9693]*kernel[2]+tmp[9791]*kernel[3]+tmp[9792]*kernel[4]+tmp[9793]*kernel[5]+tmp[9891]*kernel[6]+tmp[9892]*kernel[7]+tmp[9893]*kernel[8];
				ans[9793]<=tmp[9692]*kernel[0]+tmp[9693]*kernel[1]+tmp[9694]*kernel[2]+tmp[9792]*kernel[3]+tmp[9793]*kernel[4]+tmp[9794]*kernel[5]+tmp[9892]*kernel[6]+tmp[9893]*kernel[7]+tmp[9894]*kernel[8];
				ans[9794]<=tmp[9693]*kernel[0]+tmp[9694]*kernel[1]+tmp[9695]*kernel[2]+tmp[9793]*kernel[3]+tmp[9794]*kernel[4]+tmp[9795]*kernel[5]+tmp[9893]*kernel[6]+tmp[9894]*kernel[7]+tmp[9895]*kernel[8];
				ans[9795]<=tmp[9694]*kernel[0]+tmp[9695]*kernel[1]+tmp[9696]*kernel[2]+tmp[9794]*kernel[3]+tmp[9795]*kernel[4]+tmp[9796]*kernel[5]+tmp[9894]*kernel[6]+tmp[9895]*kernel[7]+tmp[9896]*kernel[8];
				ans[9796]<=tmp[9695]*kernel[0]+tmp[9696]*kernel[1]+tmp[9697]*kernel[2]+tmp[9795]*kernel[3]+tmp[9796]*kernel[4]+tmp[9797]*kernel[5]+tmp[9895]*kernel[6]+tmp[9896]*kernel[7]+tmp[9897]*kernel[8];
				ans[9797]<=tmp[9696]*kernel[0]+tmp[9697]*kernel[1]+tmp[9698]*kernel[2]+tmp[9796]*kernel[3]+tmp[9797]*kernel[4]+tmp[9798]*kernel[5]+tmp[9896]*kernel[6]+tmp[9897]*kernel[7]+tmp[9898]*kernel[8];
				ans[9798]<=tmp[9697]*kernel[0]+tmp[9698]*kernel[1]+tmp[9699]*kernel[2]+tmp[9797]*kernel[3]+tmp[9798]*kernel[4]+tmp[9799]*kernel[5]+tmp[9897]*kernel[6]+tmp[9898]*kernel[7]+tmp[9899]*kernel[8];
				ans[9799]<=tmp[9698]*kernel[0]+tmp[9699]*kernel[1]+tmp[9798]*kernel[3]+tmp[9799]*kernel[4]+tmp[9898]*kernel[6]+tmp[9899]*kernel[7];
				ans[9800]<=tmp[9700]*kernel[1]+tmp[9701]*kernel[2]+tmp[9800]*kernel[4]+tmp[9801]*kernel[5]+tmp[9900]*kernel[7]+tmp[9901]*kernel[8];
				ans[9801]<=tmp[9700]*kernel[0]+tmp[9701]*kernel[1]+tmp[9702]*kernel[2]+tmp[9800]*kernel[3]+tmp[9801]*kernel[4]+tmp[9802]*kernel[5]+tmp[9900]*kernel[6]+tmp[9901]*kernel[7]+tmp[9902]*kernel[8];
				ans[9802]<=tmp[9701]*kernel[0]+tmp[9702]*kernel[1]+tmp[9703]*kernel[2]+tmp[9801]*kernel[3]+tmp[9802]*kernel[4]+tmp[9803]*kernel[5]+tmp[9901]*kernel[6]+tmp[9902]*kernel[7]+tmp[9903]*kernel[8];
				ans[9803]<=tmp[9702]*kernel[0]+tmp[9703]*kernel[1]+tmp[9704]*kernel[2]+tmp[9802]*kernel[3]+tmp[9803]*kernel[4]+tmp[9804]*kernel[5]+tmp[9902]*kernel[6]+tmp[9903]*kernel[7]+tmp[9904]*kernel[8];
				ans[9804]<=tmp[9703]*kernel[0]+tmp[9704]*kernel[1]+tmp[9705]*kernel[2]+tmp[9803]*kernel[3]+tmp[9804]*kernel[4]+tmp[9805]*kernel[5]+tmp[9903]*kernel[6]+tmp[9904]*kernel[7]+tmp[9905]*kernel[8];
				ans[9805]<=tmp[9704]*kernel[0]+tmp[9705]*kernel[1]+tmp[9706]*kernel[2]+tmp[9804]*kernel[3]+tmp[9805]*kernel[4]+tmp[9806]*kernel[5]+tmp[9904]*kernel[6]+tmp[9905]*kernel[7]+tmp[9906]*kernel[8];
				ans[9806]<=tmp[9705]*kernel[0]+tmp[9706]*kernel[1]+tmp[9707]*kernel[2]+tmp[9805]*kernel[3]+tmp[9806]*kernel[4]+tmp[9807]*kernel[5]+tmp[9905]*kernel[6]+tmp[9906]*kernel[7]+tmp[9907]*kernel[8];
				ans[9807]<=tmp[9706]*kernel[0]+tmp[9707]*kernel[1]+tmp[9708]*kernel[2]+tmp[9806]*kernel[3]+tmp[9807]*kernel[4]+tmp[9808]*kernel[5]+tmp[9906]*kernel[6]+tmp[9907]*kernel[7]+tmp[9908]*kernel[8];
				ans[9808]<=tmp[9707]*kernel[0]+tmp[9708]*kernel[1]+tmp[9709]*kernel[2]+tmp[9807]*kernel[3]+tmp[9808]*kernel[4]+tmp[9809]*kernel[5]+tmp[9907]*kernel[6]+tmp[9908]*kernel[7]+tmp[9909]*kernel[8];
				ans[9809]<=tmp[9708]*kernel[0]+tmp[9709]*kernel[1]+tmp[9710]*kernel[2]+tmp[9808]*kernel[3]+tmp[9809]*kernel[4]+tmp[9810]*kernel[5]+tmp[9908]*kernel[6]+tmp[9909]*kernel[7]+tmp[9910]*kernel[8];
				ans[9810]<=tmp[9709]*kernel[0]+tmp[9710]*kernel[1]+tmp[9711]*kernel[2]+tmp[9809]*kernel[3]+tmp[9810]*kernel[4]+tmp[9811]*kernel[5]+tmp[9909]*kernel[6]+tmp[9910]*kernel[7]+tmp[9911]*kernel[8];
				ans[9811]<=tmp[9710]*kernel[0]+tmp[9711]*kernel[1]+tmp[9712]*kernel[2]+tmp[9810]*kernel[3]+tmp[9811]*kernel[4]+tmp[9812]*kernel[5]+tmp[9910]*kernel[6]+tmp[9911]*kernel[7]+tmp[9912]*kernel[8];
				ans[9812]<=tmp[9711]*kernel[0]+tmp[9712]*kernel[1]+tmp[9713]*kernel[2]+tmp[9811]*kernel[3]+tmp[9812]*kernel[4]+tmp[9813]*kernel[5]+tmp[9911]*kernel[6]+tmp[9912]*kernel[7]+tmp[9913]*kernel[8];
				ans[9813]<=tmp[9712]*kernel[0]+tmp[9713]*kernel[1]+tmp[9714]*kernel[2]+tmp[9812]*kernel[3]+tmp[9813]*kernel[4]+tmp[9814]*kernel[5]+tmp[9912]*kernel[6]+tmp[9913]*kernel[7]+tmp[9914]*kernel[8];
				ans[9814]<=tmp[9713]*kernel[0]+tmp[9714]*kernel[1]+tmp[9715]*kernel[2]+tmp[9813]*kernel[3]+tmp[9814]*kernel[4]+tmp[9815]*kernel[5]+tmp[9913]*kernel[6]+tmp[9914]*kernel[7]+tmp[9915]*kernel[8];
				ans[9815]<=tmp[9714]*kernel[0]+tmp[9715]*kernel[1]+tmp[9716]*kernel[2]+tmp[9814]*kernel[3]+tmp[9815]*kernel[4]+tmp[9816]*kernel[5]+tmp[9914]*kernel[6]+tmp[9915]*kernel[7]+tmp[9916]*kernel[8];
				ans[9816]<=tmp[9715]*kernel[0]+tmp[9716]*kernel[1]+tmp[9717]*kernel[2]+tmp[9815]*kernel[3]+tmp[9816]*kernel[4]+tmp[9817]*kernel[5]+tmp[9915]*kernel[6]+tmp[9916]*kernel[7]+tmp[9917]*kernel[8];
				ans[9817]<=tmp[9716]*kernel[0]+tmp[9717]*kernel[1]+tmp[9718]*kernel[2]+tmp[9816]*kernel[3]+tmp[9817]*kernel[4]+tmp[9818]*kernel[5]+tmp[9916]*kernel[6]+tmp[9917]*kernel[7]+tmp[9918]*kernel[8];
				ans[9818]<=tmp[9717]*kernel[0]+tmp[9718]*kernel[1]+tmp[9719]*kernel[2]+tmp[9817]*kernel[3]+tmp[9818]*kernel[4]+tmp[9819]*kernel[5]+tmp[9917]*kernel[6]+tmp[9918]*kernel[7]+tmp[9919]*kernel[8];
				ans[9819]<=tmp[9718]*kernel[0]+tmp[9719]*kernel[1]+tmp[9720]*kernel[2]+tmp[9818]*kernel[3]+tmp[9819]*kernel[4]+tmp[9820]*kernel[5]+tmp[9918]*kernel[6]+tmp[9919]*kernel[7]+tmp[9920]*kernel[8];
				ans[9820]<=tmp[9719]*kernel[0]+tmp[9720]*kernel[1]+tmp[9721]*kernel[2]+tmp[9819]*kernel[3]+tmp[9820]*kernel[4]+tmp[9821]*kernel[5]+tmp[9919]*kernel[6]+tmp[9920]*kernel[7]+tmp[9921]*kernel[8];
				ans[9821]<=tmp[9720]*kernel[0]+tmp[9721]*kernel[1]+tmp[9722]*kernel[2]+tmp[9820]*kernel[3]+tmp[9821]*kernel[4]+tmp[9822]*kernel[5]+tmp[9920]*kernel[6]+tmp[9921]*kernel[7]+tmp[9922]*kernel[8];
				ans[9822]<=tmp[9721]*kernel[0]+tmp[9722]*kernel[1]+tmp[9723]*kernel[2]+tmp[9821]*kernel[3]+tmp[9822]*kernel[4]+tmp[9823]*kernel[5]+tmp[9921]*kernel[6]+tmp[9922]*kernel[7]+tmp[9923]*kernel[8];
				ans[9823]<=tmp[9722]*kernel[0]+tmp[9723]*kernel[1]+tmp[9724]*kernel[2]+tmp[9822]*kernel[3]+tmp[9823]*kernel[4]+tmp[9824]*kernel[5]+tmp[9922]*kernel[6]+tmp[9923]*kernel[7]+tmp[9924]*kernel[8];
				ans[9824]<=tmp[9723]*kernel[0]+tmp[9724]*kernel[1]+tmp[9725]*kernel[2]+tmp[9823]*kernel[3]+tmp[9824]*kernel[4]+tmp[9825]*kernel[5]+tmp[9923]*kernel[6]+tmp[9924]*kernel[7]+tmp[9925]*kernel[8];
				ans[9825]<=tmp[9724]*kernel[0]+tmp[9725]*kernel[1]+tmp[9726]*kernel[2]+tmp[9824]*kernel[3]+tmp[9825]*kernel[4]+tmp[9826]*kernel[5]+tmp[9924]*kernel[6]+tmp[9925]*kernel[7]+tmp[9926]*kernel[8];
				ans[9826]<=tmp[9725]*kernel[0]+tmp[9726]*kernel[1]+tmp[9727]*kernel[2]+tmp[9825]*kernel[3]+tmp[9826]*kernel[4]+tmp[9827]*kernel[5]+tmp[9925]*kernel[6]+tmp[9926]*kernel[7]+tmp[9927]*kernel[8];
				ans[9827]<=tmp[9726]*kernel[0]+tmp[9727]*kernel[1]+tmp[9728]*kernel[2]+tmp[9826]*kernel[3]+tmp[9827]*kernel[4]+tmp[9828]*kernel[5]+tmp[9926]*kernel[6]+tmp[9927]*kernel[7]+tmp[9928]*kernel[8];
				ans[9828]<=tmp[9727]*kernel[0]+tmp[9728]*kernel[1]+tmp[9729]*kernel[2]+tmp[9827]*kernel[3]+tmp[9828]*kernel[4]+tmp[9829]*kernel[5]+tmp[9927]*kernel[6]+tmp[9928]*kernel[7]+tmp[9929]*kernel[8];
				ans[9829]<=tmp[9728]*kernel[0]+tmp[9729]*kernel[1]+tmp[9730]*kernel[2]+tmp[9828]*kernel[3]+tmp[9829]*kernel[4]+tmp[9830]*kernel[5]+tmp[9928]*kernel[6]+tmp[9929]*kernel[7]+tmp[9930]*kernel[8];
				ans[9830]<=tmp[9729]*kernel[0]+tmp[9730]*kernel[1]+tmp[9731]*kernel[2]+tmp[9829]*kernel[3]+tmp[9830]*kernel[4]+tmp[9831]*kernel[5]+tmp[9929]*kernel[6]+tmp[9930]*kernel[7]+tmp[9931]*kernel[8];
				ans[9831]<=tmp[9730]*kernel[0]+tmp[9731]*kernel[1]+tmp[9732]*kernel[2]+tmp[9830]*kernel[3]+tmp[9831]*kernel[4]+tmp[9832]*kernel[5]+tmp[9930]*kernel[6]+tmp[9931]*kernel[7]+tmp[9932]*kernel[8];
				ans[9832]<=tmp[9731]*kernel[0]+tmp[9732]*kernel[1]+tmp[9733]*kernel[2]+tmp[9831]*kernel[3]+tmp[9832]*kernel[4]+tmp[9833]*kernel[5]+tmp[9931]*kernel[6]+tmp[9932]*kernel[7]+tmp[9933]*kernel[8];
				ans[9833]<=tmp[9732]*kernel[0]+tmp[9733]*kernel[1]+tmp[9734]*kernel[2]+tmp[9832]*kernel[3]+tmp[9833]*kernel[4]+tmp[9834]*kernel[5]+tmp[9932]*kernel[6]+tmp[9933]*kernel[7]+tmp[9934]*kernel[8];
				ans[9834]<=tmp[9733]*kernel[0]+tmp[9734]*kernel[1]+tmp[9735]*kernel[2]+tmp[9833]*kernel[3]+tmp[9834]*kernel[4]+tmp[9835]*kernel[5]+tmp[9933]*kernel[6]+tmp[9934]*kernel[7]+tmp[9935]*kernel[8];
				ans[9835]<=tmp[9734]*kernel[0]+tmp[9735]*kernel[1]+tmp[9736]*kernel[2]+tmp[9834]*kernel[3]+tmp[9835]*kernel[4]+tmp[9836]*kernel[5]+tmp[9934]*kernel[6]+tmp[9935]*kernel[7]+tmp[9936]*kernel[8];
				ans[9836]<=tmp[9735]*kernel[0]+tmp[9736]*kernel[1]+tmp[9737]*kernel[2]+tmp[9835]*kernel[3]+tmp[9836]*kernel[4]+tmp[9837]*kernel[5]+tmp[9935]*kernel[6]+tmp[9936]*kernel[7]+tmp[9937]*kernel[8];
				ans[9837]<=tmp[9736]*kernel[0]+tmp[9737]*kernel[1]+tmp[9738]*kernel[2]+tmp[9836]*kernel[3]+tmp[9837]*kernel[4]+tmp[9838]*kernel[5]+tmp[9936]*kernel[6]+tmp[9937]*kernel[7]+tmp[9938]*kernel[8];
				ans[9838]<=tmp[9737]*kernel[0]+tmp[9738]*kernel[1]+tmp[9739]*kernel[2]+tmp[9837]*kernel[3]+tmp[9838]*kernel[4]+tmp[9839]*kernel[5]+tmp[9937]*kernel[6]+tmp[9938]*kernel[7]+tmp[9939]*kernel[8];
				ans[9839]<=tmp[9738]*kernel[0]+tmp[9739]*kernel[1]+tmp[9740]*kernel[2]+tmp[9838]*kernel[3]+tmp[9839]*kernel[4]+tmp[9840]*kernel[5]+tmp[9938]*kernel[6]+tmp[9939]*kernel[7]+tmp[9940]*kernel[8];
				ans[9840]<=tmp[9739]*kernel[0]+tmp[9740]*kernel[1]+tmp[9741]*kernel[2]+tmp[9839]*kernel[3]+tmp[9840]*kernel[4]+tmp[9841]*kernel[5]+tmp[9939]*kernel[6]+tmp[9940]*kernel[7]+tmp[9941]*kernel[8];
				ans[9841]<=tmp[9740]*kernel[0]+tmp[9741]*kernel[1]+tmp[9742]*kernel[2]+tmp[9840]*kernel[3]+tmp[9841]*kernel[4]+tmp[9842]*kernel[5]+tmp[9940]*kernel[6]+tmp[9941]*kernel[7]+tmp[9942]*kernel[8];
				ans[9842]<=tmp[9741]*kernel[0]+tmp[9742]*kernel[1]+tmp[9743]*kernel[2]+tmp[9841]*kernel[3]+tmp[9842]*kernel[4]+tmp[9843]*kernel[5]+tmp[9941]*kernel[6]+tmp[9942]*kernel[7]+tmp[9943]*kernel[8];
				ans[9843]<=tmp[9742]*kernel[0]+tmp[9743]*kernel[1]+tmp[9744]*kernel[2]+tmp[9842]*kernel[3]+tmp[9843]*kernel[4]+tmp[9844]*kernel[5]+tmp[9942]*kernel[6]+tmp[9943]*kernel[7]+tmp[9944]*kernel[8];
				ans[9844]<=tmp[9743]*kernel[0]+tmp[9744]*kernel[1]+tmp[9745]*kernel[2]+tmp[9843]*kernel[3]+tmp[9844]*kernel[4]+tmp[9845]*kernel[5]+tmp[9943]*kernel[6]+tmp[9944]*kernel[7]+tmp[9945]*kernel[8];
				ans[9845]<=tmp[9744]*kernel[0]+tmp[9745]*kernel[1]+tmp[9746]*kernel[2]+tmp[9844]*kernel[3]+tmp[9845]*kernel[4]+tmp[9846]*kernel[5]+tmp[9944]*kernel[6]+tmp[9945]*kernel[7]+tmp[9946]*kernel[8];
				ans[9846]<=tmp[9745]*kernel[0]+tmp[9746]*kernel[1]+tmp[9747]*kernel[2]+tmp[9845]*kernel[3]+tmp[9846]*kernel[4]+tmp[9847]*kernel[5]+tmp[9945]*kernel[6]+tmp[9946]*kernel[7]+tmp[9947]*kernel[8];
				ans[9847]<=tmp[9746]*kernel[0]+tmp[9747]*kernel[1]+tmp[9748]*kernel[2]+tmp[9846]*kernel[3]+tmp[9847]*kernel[4]+tmp[9848]*kernel[5]+tmp[9946]*kernel[6]+tmp[9947]*kernel[7]+tmp[9948]*kernel[8];
				ans[9848]<=tmp[9747]*kernel[0]+tmp[9748]*kernel[1]+tmp[9749]*kernel[2]+tmp[9847]*kernel[3]+tmp[9848]*kernel[4]+tmp[9849]*kernel[5]+tmp[9947]*kernel[6]+tmp[9948]*kernel[7]+tmp[9949]*kernel[8];
				ans[9849]<=tmp[9748]*kernel[0]+tmp[9749]*kernel[1]+tmp[9750]*kernel[2]+tmp[9848]*kernel[3]+tmp[9849]*kernel[4]+tmp[9850]*kernel[5]+tmp[9948]*kernel[6]+tmp[9949]*kernel[7]+tmp[9950]*kernel[8];
				ans[9850]<=tmp[9749]*kernel[0]+tmp[9750]*kernel[1]+tmp[9751]*kernel[2]+tmp[9849]*kernel[3]+tmp[9850]*kernel[4]+tmp[9851]*kernel[5]+tmp[9949]*kernel[6]+tmp[9950]*kernel[7]+tmp[9951]*kernel[8];
				ans[9851]<=tmp[9750]*kernel[0]+tmp[9751]*kernel[1]+tmp[9752]*kernel[2]+tmp[9850]*kernel[3]+tmp[9851]*kernel[4]+tmp[9852]*kernel[5]+tmp[9950]*kernel[6]+tmp[9951]*kernel[7]+tmp[9952]*kernel[8];
				ans[9852]<=tmp[9751]*kernel[0]+tmp[9752]*kernel[1]+tmp[9753]*kernel[2]+tmp[9851]*kernel[3]+tmp[9852]*kernel[4]+tmp[9853]*kernel[5]+tmp[9951]*kernel[6]+tmp[9952]*kernel[7]+tmp[9953]*kernel[8];
				ans[9853]<=tmp[9752]*kernel[0]+tmp[9753]*kernel[1]+tmp[9754]*kernel[2]+tmp[9852]*kernel[3]+tmp[9853]*kernel[4]+tmp[9854]*kernel[5]+tmp[9952]*kernel[6]+tmp[9953]*kernel[7]+tmp[9954]*kernel[8];
				ans[9854]<=tmp[9753]*kernel[0]+tmp[9754]*kernel[1]+tmp[9755]*kernel[2]+tmp[9853]*kernel[3]+tmp[9854]*kernel[4]+tmp[9855]*kernel[5]+tmp[9953]*kernel[6]+tmp[9954]*kernel[7]+tmp[9955]*kernel[8];
				ans[9855]<=tmp[9754]*kernel[0]+tmp[9755]*kernel[1]+tmp[9756]*kernel[2]+tmp[9854]*kernel[3]+tmp[9855]*kernel[4]+tmp[9856]*kernel[5]+tmp[9954]*kernel[6]+tmp[9955]*kernel[7]+tmp[9956]*kernel[8];
				ans[9856]<=tmp[9755]*kernel[0]+tmp[9756]*kernel[1]+tmp[9757]*kernel[2]+tmp[9855]*kernel[3]+tmp[9856]*kernel[4]+tmp[9857]*kernel[5]+tmp[9955]*kernel[6]+tmp[9956]*kernel[7]+tmp[9957]*kernel[8];
				ans[9857]<=tmp[9756]*kernel[0]+tmp[9757]*kernel[1]+tmp[9758]*kernel[2]+tmp[9856]*kernel[3]+tmp[9857]*kernel[4]+tmp[9858]*kernel[5]+tmp[9956]*kernel[6]+tmp[9957]*kernel[7]+tmp[9958]*kernel[8];
				ans[9858]<=tmp[9757]*kernel[0]+tmp[9758]*kernel[1]+tmp[9759]*kernel[2]+tmp[9857]*kernel[3]+tmp[9858]*kernel[4]+tmp[9859]*kernel[5]+tmp[9957]*kernel[6]+tmp[9958]*kernel[7]+tmp[9959]*kernel[8];
				ans[9859]<=tmp[9758]*kernel[0]+tmp[9759]*kernel[1]+tmp[9760]*kernel[2]+tmp[9858]*kernel[3]+tmp[9859]*kernel[4]+tmp[9860]*kernel[5]+tmp[9958]*kernel[6]+tmp[9959]*kernel[7]+tmp[9960]*kernel[8];
				ans[9860]<=tmp[9759]*kernel[0]+tmp[9760]*kernel[1]+tmp[9761]*kernel[2]+tmp[9859]*kernel[3]+tmp[9860]*kernel[4]+tmp[9861]*kernel[5]+tmp[9959]*kernel[6]+tmp[9960]*kernel[7]+tmp[9961]*kernel[8];
				ans[9861]<=tmp[9760]*kernel[0]+tmp[9761]*kernel[1]+tmp[9762]*kernel[2]+tmp[9860]*kernel[3]+tmp[9861]*kernel[4]+tmp[9862]*kernel[5]+tmp[9960]*kernel[6]+tmp[9961]*kernel[7]+tmp[9962]*kernel[8];
				ans[9862]<=tmp[9761]*kernel[0]+tmp[9762]*kernel[1]+tmp[9763]*kernel[2]+tmp[9861]*kernel[3]+tmp[9862]*kernel[4]+tmp[9863]*kernel[5]+tmp[9961]*kernel[6]+tmp[9962]*kernel[7]+tmp[9963]*kernel[8];
				ans[9863]<=tmp[9762]*kernel[0]+tmp[9763]*kernel[1]+tmp[9764]*kernel[2]+tmp[9862]*kernel[3]+tmp[9863]*kernel[4]+tmp[9864]*kernel[5]+tmp[9962]*kernel[6]+tmp[9963]*kernel[7]+tmp[9964]*kernel[8];
				ans[9864]<=tmp[9763]*kernel[0]+tmp[9764]*kernel[1]+tmp[9765]*kernel[2]+tmp[9863]*kernel[3]+tmp[9864]*kernel[4]+tmp[9865]*kernel[5]+tmp[9963]*kernel[6]+tmp[9964]*kernel[7]+tmp[9965]*kernel[8];
				ans[9865]<=tmp[9764]*kernel[0]+tmp[9765]*kernel[1]+tmp[9766]*kernel[2]+tmp[9864]*kernel[3]+tmp[9865]*kernel[4]+tmp[9866]*kernel[5]+tmp[9964]*kernel[6]+tmp[9965]*kernel[7]+tmp[9966]*kernel[8];
				ans[9866]<=tmp[9765]*kernel[0]+tmp[9766]*kernel[1]+tmp[9767]*kernel[2]+tmp[9865]*kernel[3]+tmp[9866]*kernel[4]+tmp[9867]*kernel[5]+tmp[9965]*kernel[6]+tmp[9966]*kernel[7]+tmp[9967]*kernel[8];
				ans[9867]<=tmp[9766]*kernel[0]+tmp[9767]*kernel[1]+tmp[9768]*kernel[2]+tmp[9866]*kernel[3]+tmp[9867]*kernel[4]+tmp[9868]*kernel[5]+tmp[9966]*kernel[6]+tmp[9967]*kernel[7]+tmp[9968]*kernel[8];
				ans[9868]<=tmp[9767]*kernel[0]+tmp[9768]*kernel[1]+tmp[9769]*kernel[2]+tmp[9867]*kernel[3]+tmp[9868]*kernel[4]+tmp[9869]*kernel[5]+tmp[9967]*kernel[6]+tmp[9968]*kernel[7]+tmp[9969]*kernel[8];
				ans[9869]<=tmp[9768]*kernel[0]+tmp[9769]*kernel[1]+tmp[9770]*kernel[2]+tmp[9868]*kernel[3]+tmp[9869]*kernel[4]+tmp[9870]*kernel[5]+tmp[9968]*kernel[6]+tmp[9969]*kernel[7]+tmp[9970]*kernel[8];
				ans[9870]<=tmp[9769]*kernel[0]+tmp[9770]*kernel[1]+tmp[9771]*kernel[2]+tmp[9869]*kernel[3]+tmp[9870]*kernel[4]+tmp[9871]*kernel[5]+tmp[9969]*kernel[6]+tmp[9970]*kernel[7]+tmp[9971]*kernel[8];
				ans[9871]<=tmp[9770]*kernel[0]+tmp[9771]*kernel[1]+tmp[9772]*kernel[2]+tmp[9870]*kernel[3]+tmp[9871]*kernel[4]+tmp[9872]*kernel[5]+tmp[9970]*kernel[6]+tmp[9971]*kernel[7]+tmp[9972]*kernel[8];
				ans[9872]<=tmp[9771]*kernel[0]+tmp[9772]*kernel[1]+tmp[9773]*kernel[2]+tmp[9871]*kernel[3]+tmp[9872]*kernel[4]+tmp[9873]*kernel[5]+tmp[9971]*kernel[6]+tmp[9972]*kernel[7]+tmp[9973]*kernel[8];
				ans[9873]<=tmp[9772]*kernel[0]+tmp[9773]*kernel[1]+tmp[9774]*kernel[2]+tmp[9872]*kernel[3]+tmp[9873]*kernel[4]+tmp[9874]*kernel[5]+tmp[9972]*kernel[6]+tmp[9973]*kernel[7]+tmp[9974]*kernel[8];
				ans[9874]<=tmp[9773]*kernel[0]+tmp[9774]*kernel[1]+tmp[9775]*kernel[2]+tmp[9873]*kernel[3]+tmp[9874]*kernel[4]+tmp[9875]*kernel[5]+tmp[9973]*kernel[6]+tmp[9974]*kernel[7]+tmp[9975]*kernel[8];
				ans[9875]<=tmp[9774]*kernel[0]+tmp[9775]*kernel[1]+tmp[9776]*kernel[2]+tmp[9874]*kernel[3]+tmp[9875]*kernel[4]+tmp[9876]*kernel[5]+tmp[9974]*kernel[6]+tmp[9975]*kernel[7]+tmp[9976]*kernel[8];
				ans[9876]<=tmp[9775]*kernel[0]+tmp[9776]*kernel[1]+tmp[9777]*kernel[2]+tmp[9875]*kernel[3]+tmp[9876]*kernel[4]+tmp[9877]*kernel[5]+tmp[9975]*kernel[6]+tmp[9976]*kernel[7]+tmp[9977]*kernel[8];
				ans[9877]<=tmp[9776]*kernel[0]+tmp[9777]*kernel[1]+tmp[9778]*kernel[2]+tmp[9876]*kernel[3]+tmp[9877]*kernel[4]+tmp[9878]*kernel[5]+tmp[9976]*kernel[6]+tmp[9977]*kernel[7]+tmp[9978]*kernel[8];
				ans[9878]<=tmp[9777]*kernel[0]+tmp[9778]*kernel[1]+tmp[9779]*kernel[2]+tmp[9877]*kernel[3]+tmp[9878]*kernel[4]+tmp[9879]*kernel[5]+tmp[9977]*kernel[6]+tmp[9978]*kernel[7]+tmp[9979]*kernel[8];
				ans[9879]<=tmp[9778]*kernel[0]+tmp[9779]*kernel[1]+tmp[9780]*kernel[2]+tmp[9878]*kernel[3]+tmp[9879]*kernel[4]+tmp[9880]*kernel[5]+tmp[9978]*kernel[6]+tmp[9979]*kernel[7]+tmp[9980]*kernel[8];
				ans[9880]<=tmp[9779]*kernel[0]+tmp[9780]*kernel[1]+tmp[9781]*kernel[2]+tmp[9879]*kernel[3]+tmp[9880]*kernel[4]+tmp[9881]*kernel[5]+tmp[9979]*kernel[6]+tmp[9980]*kernel[7]+tmp[9981]*kernel[8];
				ans[9881]<=tmp[9780]*kernel[0]+tmp[9781]*kernel[1]+tmp[9782]*kernel[2]+tmp[9880]*kernel[3]+tmp[9881]*kernel[4]+tmp[9882]*kernel[5]+tmp[9980]*kernel[6]+tmp[9981]*kernel[7]+tmp[9982]*kernel[8];
				ans[9882]<=tmp[9781]*kernel[0]+tmp[9782]*kernel[1]+tmp[9783]*kernel[2]+tmp[9881]*kernel[3]+tmp[9882]*kernel[4]+tmp[9883]*kernel[5]+tmp[9981]*kernel[6]+tmp[9982]*kernel[7]+tmp[9983]*kernel[8];
				ans[9883]<=tmp[9782]*kernel[0]+tmp[9783]*kernel[1]+tmp[9784]*kernel[2]+tmp[9882]*kernel[3]+tmp[9883]*kernel[4]+tmp[9884]*kernel[5]+tmp[9982]*kernel[6]+tmp[9983]*kernel[7]+tmp[9984]*kernel[8];
				ans[9884]<=tmp[9783]*kernel[0]+tmp[9784]*kernel[1]+tmp[9785]*kernel[2]+tmp[9883]*kernel[3]+tmp[9884]*kernel[4]+tmp[9885]*kernel[5]+tmp[9983]*kernel[6]+tmp[9984]*kernel[7]+tmp[9985]*kernel[8];
				ans[9885]<=tmp[9784]*kernel[0]+tmp[9785]*kernel[1]+tmp[9786]*kernel[2]+tmp[9884]*kernel[3]+tmp[9885]*kernel[4]+tmp[9886]*kernel[5]+tmp[9984]*kernel[6]+tmp[9985]*kernel[7]+tmp[9986]*kernel[8];
				ans[9886]<=tmp[9785]*kernel[0]+tmp[9786]*kernel[1]+tmp[9787]*kernel[2]+tmp[9885]*kernel[3]+tmp[9886]*kernel[4]+tmp[9887]*kernel[5]+tmp[9985]*kernel[6]+tmp[9986]*kernel[7]+tmp[9987]*kernel[8];
				ans[9887]<=tmp[9786]*kernel[0]+tmp[9787]*kernel[1]+tmp[9788]*kernel[2]+tmp[9886]*kernel[3]+tmp[9887]*kernel[4]+tmp[9888]*kernel[5]+tmp[9986]*kernel[6]+tmp[9987]*kernel[7]+tmp[9988]*kernel[8];
				ans[9888]<=tmp[9787]*kernel[0]+tmp[9788]*kernel[1]+tmp[9789]*kernel[2]+tmp[9887]*kernel[3]+tmp[9888]*kernel[4]+tmp[9889]*kernel[5]+tmp[9987]*kernel[6]+tmp[9988]*kernel[7]+tmp[9989]*kernel[8];
				ans[9889]<=tmp[9788]*kernel[0]+tmp[9789]*kernel[1]+tmp[9790]*kernel[2]+tmp[9888]*kernel[3]+tmp[9889]*kernel[4]+tmp[9890]*kernel[5]+tmp[9988]*kernel[6]+tmp[9989]*kernel[7]+tmp[9990]*kernel[8];
				ans[9890]<=tmp[9789]*kernel[0]+tmp[9790]*kernel[1]+tmp[9791]*kernel[2]+tmp[9889]*kernel[3]+tmp[9890]*kernel[4]+tmp[9891]*kernel[5]+tmp[9989]*kernel[6]+tmp[9990]*kernel[7]+tmp[9991]*kernel[8];
				ans[9891]<=tmp[9790]*kernel[0]+tmp[9791]*kernel[1]+tmp[9792]*kernel[2]+tmp[9890]*kernel[3]+tmp[9891]*kernel[4]+tmp[9892]*kernel[5]+tmp[9990]*kernel[6]+tmp[9991]*kernel[7]+tmp[9992]*kernel[8];
				ans[9892]<=tmp[9791]*kernel[0]+tmp[9792]*kernel[1]+tmp[9793]*kernel[2]+tmp[9891]*kernel[3]+tmp[9892]*kernel[4]+tmp[9893]*kernel[5]+tmp[9991]*kernel[6]+tmp[9992]*kernel[7]+tmp[9993]*kernel[8];
				ans[9893]<=tmp[9792]*kernel[0]+tmp[9793]*kernel[1]+tmp[9794]*kernel[2]+tmp[9892]*kernel[3]+tmp[9893]*kernel[4]+tmp[9894]*kernel[5]+tmp[9992]*kernel[6]+tmp[9993]*kernel[7]+tmp[9994]*kernel[8];
				ans[9894]<=tmp[9793]*kernel[0]+tmp[9794]*kernel[1]+tmp[9795]*kernel[2]+tmp[9893]*kernel[3]+tmp[9894]*kernel[4]+tmp[9895]*kernel[5]+tmp[9993]*kernel[6]+tmp[9994]*kernel[7]+tmp[9995]*kernel[8];
				ans[9895]<=tmp[9794]*kernel[0]+tmp[9795]*kernel[1]+tmp[9796]*kernel[2]+tmp[9894]*kernel[3]+tmp[9895]*kernel[4]+tmp[9896]*kernel[5]+tmp[9994]*kernel[6]+tmp[9995]*kernel[7]+tmp[9996]*kernel[8];
				ans[9896]<=tmp[9795]*kernel[0]+tmp[9796]*kernel[1]+tmp[9797]*kernel[2]+tmp[9895]*kernel[3]+tmp[9896]*kernel[4]+tmp[9897]*kernel[5]+tmp[9995]*kernel[6]+tmp[9996]*kernel[7]+tmp[9997]*kernel[8];
				ans[9897]<=tmp[9796]*kernel[0]+tmp[9797]*kernel[1]+tmp[9798]*kernel[2]+tmp[9896]*kernel[3]+tmp[9897]*kernel[4]+tmp[9898]*kernel[5]+tmp[9996]*kernel[6]+tmp[9997]*kernel[7]+tmp[9998]*kernel[8];
				ans[9898]<=tmp[9797]*kernel[0]+tmp[9798]*kernel[1]+tmp[9799]*kernel[2]+tmp[9897]*kernel[3]+tmp[9898]*kernel[4]+tmp[9899]*kernel[5]+tmp[9997]*kernel[6]+tmp[9998]*kernel[7]+tmp[9999]*kernel[8];
				ans[9899]<=tmp[9798]*kernel[0]+tmp[9799]*kernel[1]+tmp[9898]*kernel[3]+tmp[9899]*kernel[4]+tmp[9998]*kernel[6]+tmp[9999]*kernel[7];
				ans[9900]<=tmp[9800]*kernel[1]+tmp[9801]*kernel[2]+tmp[9900]*kernel[4]+tmp[9901]*kernel[5];
				ans[9901]<=tmp[9800]*kernel[0]+tmp[9801]*kernel[1]+tmp[9802]*kernel[2]+tmp[9900]*kernel[3]+tmp[9901]*kernel[4]+tmp[9902]*kernel[5];
				ans[9902]<=tmp[9801]*kernel[0]+tmp[9802]*kernel[1]+tmp[9803]*kernel[2]+tmp[9901]*kernel[3]+tmp[9902]*kernel[4]+tmp[9903]*kernel[5];
				ans[9903]<=tmp[9802]*kernel[0]+tmp[9803]*kernel[1]+tmp[9804]*kernel[2]+tmp[9902]*kernel[3]+tmp[9903]*kernel[4]+tmp[9904]*kernel[5];
				ans[9904]<=tmp[9803]*kernel[0]+tmp[9804]*kernel[1]+tmp[9805]*kernel[2]+tmp[9903]*kernel[3]+tmp[9904]*kernel[4]+tmp[9905]*kernel[5];
				ans[9905]<=tmp[9804]*kernel[0]+tmp[9805]*kernel[1]+tmp[9806]*kernel[2]+tmp[9904]*kernel[3]+tmp[9905]*kernel[4]+tmp[9906]*kernel[5];
				ans[9906]<=tmp[9805]*kernel[0]+tmp[9806]*kernel[1]+tmp[9807]*kernel[2]+tmp[9905]*kernel[3]+tmp[9906]*kernel[4]+tmp[9907]*kernel[5];
				ans[9907]<=tmp[9806]*kernel[0]+tmp[9807]*kernel[1]+tmp[9808]*kernel[2]+tmp[9906]*kernel[3]+tmp[9907]*kernel[4]+tmp[9908]*kernel[5];
				ans[9908]<=tmp[9807]*kernel[0]+tmp[9808]*kernel[1]+tmp[9809]*kernel[2]+tmp[9907]*kernel[3]+tmp[9908]*kernel[4]+tmp[9909]*kernel[5];
				ans[9909]<=tmp[9808]*kernel[0]+tmp[9809]*kernel[1]+tmp[9810]*kernel[2]+tmp[9908]*kernel[3]+tmp[9909]*kernel[4]+tmp[9910]*kernel[5];
				ans[9910]<=tmp[9809]*kernel[0]+tmp[9810]*kernel[1]+tmp[9811]*kernel[2]+tmp[9909]*kernel[3]+tmp[9910]*kernel[4]+tmp[9911]*kernel[5];
				ans[9911]<=tmp[9810]*kernel[0]+tmp[9811]*kernel[1]+tmp[9812]*kernel[2]+tmp[9910]*kernel[3]+tmp[9911]*kernel[4]+tmp[9912]*kernel[5];
				ans[9912]<=tmp[9811]*kernel[0]+tmp[9812]*kernel[1]+tmp[9813]*kernel[2]+tmp[9911]*kernel[3]+tmp[9912]*kernel[4]+tmp[9913]*kernel[5];
				ans[9913]<=tmp[9812]*kernel[0]+tmp[9813]*kernel[1]+tmp[9814]*kernel[2]+tmp[9912]*kernel[3]+tmp[9913]*kernel[4]+tmp[9914]*kernel[5];
				ans[9914]<=tmp[9813]*kernel[0]+tmp[9814]*kernel[1]+tmp[9815]*kernel[2]+tmp[9913]*kernel[3]+tmp[9914]*kernel[4]+tmp[9915]*kernel[5];
				ans[9915]<=tmp[9814]*kernel[0]+tmp[9815]*kernel[1]+tmp[9816]*kernel[2]+tmp[9914]*kernel[3]+tmp[9915]*kernel[4]+tmp[9916]*kernel[5];
				ans[9916]<=tmp[9815]*kernel[0]+tmp[9816]*kernel[1]+tmp[9817]*kernel[2]+tmp[9915]*kernel[3]+tmp[9916]*kernel[4]+tmp[9917]*kernel[5];
				ans[9917]<=tmp[9816]*kernel[0]+tmp[9817]*kernel[1]+tmp[9818]*kernel[2]+tmp[9916]*kernel[3]+tmp[9917]*kernel[4]+tmp[9918]*kernel[5];
				ans[9918]<=tmp[9817]*kernel[0]+tmp[9818]*kernel[1]+tmp[9819]*kernel[2]+tmp[9917]*kernel[3]+tmp[9918]*kernel[4]+tmp[9919]*kernel[5];
				ans[9919]<=tmp[9818]*kernel[0]+tmp[9819]*kernel[1]+tmp[9820]*kernel[2]+tmp[9918]*kernel[3]+tmp[9919]*kernel[4]+tmp[9920]*kernel[5];
				ans[9920]<=tmp[9819]*kernel[0]+tmp[9820]*kernel[1]+tmp[9821]*kernel[2]+tmp[9919]*kernel[3]+tmp[9920]*kernel[4]+tmp[9921]*kernel[5];
				ans[9921]<=tmp[9820]*kernel[0]+tmp[9821]*kernel[1]+tmp[9822]*kernel[2]+tmp[9920]*kernel[3]+tmp[9921]*kernel[4]+tmp[9922]*kernel[5];
				ans[9922]<=tmp[9821]*kernel[0]+tmp[9822]*kernel[1]+tmp[9823]*kernel[2]+tmp[9921]*kernel[3]+tmp[9922]*kernel[4]+tmp[9923]*kernel[5];
				ans[9923]<=tmp[9822]*kernel[0]+tmp[9823]*kernel[1]+tmp[9824]*kernel[2]+tmp[9922]*kernel[3]+tmp[9923]*kernel[4]+tmp[9924]*kernel[5];
				ans[9924]<=tmp[9823]*kernel[0]+tmp[9824]*kernel[1]+tmp[9825]*kernel[2]+tmp[9923]*kernel[3]+tmp[9924]*kernel[4]+tmp[9925]*kernel[5];
				ans[9925]<=tmp[9824]*kernel[0]+tmp[9825]*kernel[1]+tmp[9826]*kernel[2]+tmp[9924]*kernel[3]+tmp[9925]*kernel[4]+tmp[9926]*kernel[5];
				ans[9926]<=tmp[9825]*kernel[0]+tmp[9826]*kernel[1]+tmp[9827]*kernel[2]+tmp[9925]*kernel[3]+tmp[9926]*kernel[4]+tmp[9927]*kernel[5];
				ans[9927]<=tmp[9826]*kernel[0]+tmp[9827]*kernel[1]+tmp[9828]*kernel[2]+tmp[9926]*kernel[3]+tmp[9927]*kernel[4]+tmp[9928]*kernel[5];
				ans[9928]<=tmp[9827]*kernel[0]+tmp[9828]*kernel[1]+tmp[9829]*kernel[2]+tmp[9927]*kernel[3]+tmp[9928]*kernel[4]+tmp[9929]*kernel[5];
				ans[9929]<=tmp[9828]*kernel[0]+tmp[9829]*kernel[1]+tmp[9830]*kernel[2]+tmp[9928]*kernel[3]+tmp[9929]*kernel[4]+tmp[9930]*kernel[5];
				ans[9930]<=tmp[9829]*kernel[0]+tmp[9830]*kernel[1]+tmp[9831]*kernel[2]+tmp[9929]*kernel[3]+tmp[9930]*kernel[4]+tmp[9931]*kernel[5];
				ans[9931]<=tmp[9830]*kernel[0]+tmp[9831]*kernel[1]+tmp[9832]*kernel[2]+tmp[9930]*kernel[3]+tmp[9931]*kernel[4]+tmp[9932]*kernel[5];
				ans[9932]<=tmp[9831]*kernel[0]+tmp[9832]*kernel[1]+tmp[9833]*kernel[2]+tmp[9931]*kernel[3]+tmp[9932]*kernel[4]+tmp[9933]*kernel[5];
				ans[9933]<=tmp[9832]*kernel[0]+tmp[9833]*kernel[1]+tmp[9834]*kernel[2]+tmp[9932]*kernel[3]+tmp[9933]*kernel[4]+tmp[9934]*kernel[5];
				ans[9934]<=tmp[9833]*kernel[0]+tmp[9834]*kernel[1]+tmp[9835]*kernel[2]+tmp[9933]*kernel[3]+tmp[9934]*kernel[4]+tmp[9935]*kernel[5];
				ans[9935]<=tmp[9834]*kernel[0]+tmp[9835]*kernel[1]+tmp[9836]*kernel[2]+tmp[9934]*kernel[3]+tmp[9935]*kernel[4]+tmp[9936]*kernel[5];
				ans[9936]<=tmp[9835]*kernel[0]+tmp[9836]*kernel[1]+tmp[9837]*kernel[2]+tmp[9935]*kernel[3]+tmp[9936]*kernel[4]+tmp[9937]*kernel[5];
				ans[9937]<=tmp[9836]*kernel[0]+tmp[9837]*kernel[1]+tmp[9838]*kernel[2]+tmp[9936]*kernel[3]+tmp[9937]*kernel[4]+tmp[9938]*kernel[5];
				ans[9938]<=tmp[9837]*kernel[0]+tmp[9838]*kernel[1]+tmp[9839]*kernel[2]+tmp[9937]*kernel[3]+tmp[9938]*kernel[4]+tmp[9939]*kernel[5];
				ans[9939]<=tmp[9838]*kernel[0]+tmp[9839]*kernel[1]+tmp[9840]*kernel[2]+tmp[9938]*kernel[3]+tmp[9939]*kernel[4]+tmp[9940]*kernel[5];
				ans[9940]<=tmp[9839]*kernel[0]+tmp[9840]*kernel[1]+tmp[9841]*kernel[2]+tmp[9939]*kernel[3]+tmp[9940]*kernel[4]+tmp[9941]*kernel[5];
				ans[9941]<=tmp[9840]*kernel[0]+tmp[9841]*kernel[1]+tmp[9842]*kernel[2]+tmp[9940]*kernel[3]+tmp[9941]*kernel[4]+tmp[9942]*kernel[5];
				ans[9942]<=tmp[9841]*kernel[0]+tmp[9842]*kernel[1]+tmp[9843]*kernel[2]+tmp[9941]*kernel[3]+tmp[9942]*kernel[4]+tmp[9943]*kernel[5];
				ans[9943]<=tmp[9842]*kernel[0]+tmp[9843]*kernel[1]+tmp[9844]*kernel[2]+tmp[9942]*kernel[3]+tmp[9943]*kernel[4]+tmp[9944]*kernel[5];
				ans[9944]<=tmp[9843]*kernel[0]+tmp[9844]*kernel[1]+tmp[9845]*kernel[2]+tmp[9943]*kernel[3]+tmp[9944]*kernel[4]+tmp[9945]*kernel[5];
				ans[9945]<=tmp[9844]*kernel[0]+tmp[9845]*kernel[1]+tmp[9846]*kernel[2]+tmp[9944]*kernel[3]+tmp[9945]*kernel[4]+tmp[9946]*kernel[5];
				ans[9946]<=tmp[9845]*kernel[0]+tmp[9846]*kernel[1]+tmp[9847]*kernel[2]+tmp[9945]*kernel[3]+tmp[9946]*kernel[4]+tmp[9947]*kernel[5];
				ans[9947]<=tmp[9846]*kernel[0]+tmp[9847]*kernel[1]+tmp[9848]*kernel[2]+tmp[9946]*kernel[3]+tmp[9947]*kernel[4]+tmp[9948]*kernel[5];
				ans[9948]<=tmp[9847]*kernel[0]+tmp[9848]*kernel[1]+tmp[9849]*kernel[2]+tmp[9947]*kernel[3]+tmp[9948]*kernel[4]+tmp[9949]*kernel[5];
				ans[9949]<=tmp[9848]*kernel[0]+tmp[9849]*kernel[1]+tmp[9850]*kernel[2]+tmp[9948]*kernel[3]+tmp[9949]*kernel[4]+tmp[9950]*kernel[5];
				ans[9950]<=tmp[9849]*kernel[0]+tmp[9850]*kernel[1]+tmp[9851]*kernel[2]+tmp[9949]*kernel[3]+tmp[9950]*kernel[4]+tmp[9951]*kernel[5];
				ans[9951]<=tmp[9850]*kernel[0]+tmp[9851]*kernel[1]+tmp[9852]*kernel[2]+tmp[9950]*kernel[3]+tmp[9951]*kernel[4]+tmp[9952]*kernel[5];
				ans[9952]<=tmp[9851]*kernel[0]+tmp[9852]*kernel[1]+tmp[9853]*kernel[2]+tmp[9951]*kernel[3]+tmp[9952]*kernel[4]+tmp[9953]*kernel[5];
				ans[9953]<=tmp[9852]*kernel[0]+tmp[9853]*kernel[1]+tmp[9854]*kernel[2]+tmp[9952]*kernel[3]+tmp[9953]*kernel[4]+tmp[9954]*kernel[5];
				ans[9954]<=tmp[9853]*kernel[0]+tmp[9854]*kernel[1]+tmp[9855]*kernel[2]+tmp[9953]*kernel[3]+tmp[9954]*kernel[4]+tmp[9955]*kernel[5];
				ans[9955]<=tmp[9854]*kernel[0]+tmp[9855]*kernel[1]+tmp[9856]*kernel[2]+tmp[9954]*kernel[3]+tmp[9955]*kernel[4]+tmp[9956]*kernel[5];
				ans[9956]<=tmp[9855]*kernel[0]+tmp[9856]*kernel[1]+tmp[9857]*kernel[2]+tmp[9955]*kernel[3]+tmp[9956]*kernel[4]+tmp[9957]*kernel[5];
				ans[9957]<=tmp[9856]*kernel[0]+tmp[9857]*kernel[1]+tmp[9858]*kernel[2]+tmp[9956]*kernel[3]+tmp[9957]*kernel[4]+tmp[9958]*kernel[5];
				ans[9958]<=tmp[9857]*kernel[0]+tmp[9858]*kernel[1]+tmp[9859]*kernel[2]+tmp[9957]*kernel[3]+tmp[9958]*kernel[4]+tmp[9959]*kernel[5];
				ans[9959]<=tmp[9858]*kernel[0]+tmp[9859]*kernel[1]+tmp[9860]*kernel[2]+tmp[9958]*kernel[3]+tmp[9959]*kernel[4]+tmp[9960]*kernel[5];
				ans[9960]<=tmp[9859]*kernel[0]+tmp[9860]*kernel[1]+tmp[9861]*kernel[2]+tmp[9959]*kernel[3]+tmp[9960]*kernel[4]+tmp[9961]*kernel[5];
				ans[9961]<=tmp[9860]*kernel[0]+tmp[9861]*kernel[1]+tmp[9862]*kernel[2]+tmp[9960]*kernel[3]+tmp[9961]*kernel[4]+tmp[9962]*kernel[5];
				ans[9962]<=tmp[9861]*kernel[0]+tmp[9862]*kernel[1]+tmp[9863]*kernel[2]+tmp[9961]*kernel[3]+tmp[9962]*kernel[4]+tmp[9963]*kernel[5];
				ans[9963]<=tmp[9862]*kernel[0]+tmp[9863]*kernel[1]+tmp[9864]*kernel[2]+tmp[9962]*kernel[3]+tmp[9963]*kernel[4]+tmp[9964]*kernel[5];
				ans[9964]<=tmp[9863]*kernel[0]+tmp[9864]*kernel[1]+tmp[9865]*kernel[2]+tmp[9963]*kernel[3]+tmp[9964]*kernel[4]+tmp[9965]*kernel[5];
				ans[9965]<=tmp[9864]*kernel[0]+tmp[9865]*kernel[1]+tmp[9866]*kernel[2]+tmp[9964]*kernel[3]+tmp[9965]*kernel[4]+tmp[9966]*kernel[5];
				ans[9966]<=tmp[9865]*kernel[0]+tmp[9866]*kernel[1]+tmp[9867]*kernel[2]+tmp[9965]*kernel[3]+tmp[9966]*kernel[4]+tmp[9967]*kernel[5];
				ans[9967]<=tmp[9866]*kernel[0]+tmp[9867]*kernel[1]+tmp[9868]*kernel[2]+tmp[9966]*kernel[3]+tmp[9967]*kernel[4]+tmp[9968]*kernel[5];
				ans[9968]<=tmp[9867]*kernel[0]+tmp[9868]*kernel[1]+tmp[9869]*kernel[2]+tmp[9967]*kernel[3]+tmp[9968]*kernel[4]+tmp[9969]*kernel[5];
				ans[9969]<=tmp[9868]*kernel[0]+tmp[9869]*kernel[1]+tmp[9870]*kernel[2]+tmp[9968]*kernel[3]+tmp[9969]*kernel[4]+tmp[9970]*kernel[5];
				ans[9970]<=tmp[9869]*kernel[0]+tmp[9870]*kernel[1]+tmp[9871]*kernel[2]+tmp[9969]*kernel[3]+tmp[9970]*kernel[4]+tmp[9971]*kernel[5];
				ans[9971]<=tmp[9870]*kernel[0]+tmp[9871]*kernel[1]+tmp[9872]*kernel[2]+tmp[9970]*kernel[3]+tmp[9971]*kernel[4]+tmp[9972]*kernel[5];
				ans[9972]<=tmp[9871]*kernel[0]+tmp[9872]*kernel[1]+tmp[9873]*kernel[2]+tmp[9971]*kernel[3]+tmp[9972]*kernel[4]+tmp[9973]*kernel[5];
				ans[9973]<=tmp[9872]*kernel[0]+tmp[9873]*kernel[1]+tmp[9874]*kernel[2]+tmp[9972]*kernel[3]+tmp[9973]*kernel[4]+tmp[9974]*kernel[5];
				ans[9974]<=tmp[9873]*kernel[0]+tmp[9874]*kernel[1]+tmp[9875]*kernel[2]+tmp[9973]*kernel[3]+tmp[9974]*kernel[4]+tmp[9975]*kernel[5];
				ans[9975]<=tmp[9874]*kernel[0]+tmp[9875]*kernel[1]+tmp[9876]*kernel[2]+tmp[9974]*kernel[3]+tmp[9975]*kernel[4]+tmp[9976]*kernel[5];
				ans[9976]<=tmp[9875]*kernel[0]+tmp[9876]*kernel[1]+tmp[9877]*kernel[2]+tmp[9975]*kernel[3]+tmp[9976]*kernel[4]+tmp[9977]*kernel[5];
				ans[9977]<=tmp[9876]*kernel[0]+tmp[9877]*kernel[1]+tmp[9878]*kernel[2]+tmp[9976]*kernel[3]+tmp[9977]*kernel[4]+tmp[9978]*kernel[5];
				ans[9978]<=tmp[9877]*kernel[0]+tmp[9878]*kernel[1]+tmp[9879]*kernel[2]+tmp[9977]*kernel[3]+tmp[9978]*kernel[4]+tmp[9979]*kernel[5];
				ans[9979]<=tmp[9878]*kernel[0]+tmp[9879]*kernel[1]+tmp[9880]*kernel[2]+tmp[9978]*kernel[3]+tmp[9979]*kernel[4]+tmp[9980]*kernel[5];
				ans[9980]<=tmp[9879]*kernel[0]+tmp[9880]*kernel[1]+tmp[9881]*kernel[2]+tmp[9979]*kernel[3]+tmp[9980]*kernel[4]+tmp[9981]*kernel[5];
				ans[9981]<=tmp[9880]*kernel[0]+tmp[9881]*kernel[1]+tmp[9882]*kernel[2]+tmp[9980]*kernel[3]+tmp[9981]*kernel[4]+tmp[9982]*kernel[5];
				ans[9982]<=tmp[9881]*kernel[0]+tmp[9882]*kernel[1]+tmp[9883]*kernel[2]+tmp[9981]*kernel[3]+tmp[9982]*kernel[4]+tmp[9983]*kernel[5];
				ans[9983]<=tmp[9882]*kernel[0]+tmp[9883]*kernel[1]+tmp[9884]*kernel[2]+tmp[9982]*kernel[3]+tmp[9983]*kernel[4]+tmp[9984]*kernel[5];
				ans[9984]<=tmp[9883]*kernel[0]+tmp[9884]*kernel[1]+tmp[9885]*kernel[2]+tmp[9983]*kernel[3]+tmp[9984]*kernel[4]+tmp[9985]*kernel[5];
				ans[9985]<=tmp[9884]*kernel[0]+tmp[9885]*kernel[1]+tmp[9886]*kernel[2]+tmp[9984]*kernel[3]+tmp[9985]*kernel[4]+tmp[9986]*kernel[5];
				ans[9986]<=tmp[9885]*kernel[0]+tmp[9886]*kernel[1]+tmp[9887]*kernel[2]+tmp[9985]*kernel[3]+tmp[9986]*kernel[4]+tmp[9987]*kernel[5];
				ans[9987]<=tmp[9886]*kernel[0]+tmp[9887]*kernel[1]+tmp[9888]*kernel[2]+tmp[9986]*kernel[3]+tmp[9987]*kernel[4]+tmp[9988]*kernel[5];
				ans[9988]<=tmp[9887]*kernel[0]+tmp[9888]*kernel[1]+tmp[9889]*kernel[2]+tmp[9987]*kernel[3]+tmp[9988]*kernel[4]+tmp[9989]*kernel[5];
				ans[9989]<=tmp[9888]*kernel[0]+tmp[9889]*kernel[1]+tmp[9890]*kernel[2]+tmp[9988]*kernel[3]+tmp[9989]*kernel[4]+tmp[9990]*kernel[5];
				ans[9990]<=tmp[9889]*kernel[0]+tmp[9890]*kernel[1]+tmp[9891]*kernel[2]+tmp[9989]*kernel[3]+tmp[9990]*kernel[4]+tmp[9991]*kernel[5];
				ans[9991]<=tmp[9890]*kernel[0]+tmp[9891]*kernel[1]+tmp[9892]*kernel[2]+tmp[9990]*kernel[3]+tmp[9991]*kernel[4]+tmp[9992]*kernel[5];
				ans[9992]<=tmp[9891]*kernel[0]+tmp[9892]*kernel[1]+tmp[9893]*kernel[2]+tmp[9991]*kernel[3]+tmp[9992]*kernel[4]+tmp[9993]*kernel[5];
				ans[9993]<=tmp[9892]*kernel[0]+tmp[9893]*kernel[1]+tmp[9894]*kernel[2]+tmp[9992]*kernel[3]+tmp[9993]*kernel[4]+tmp[9994]*kernel[5];
				ans[9994]<=tmp[9893]*kernel[0]+tmp[9894]*kernel[1]+tmp[9895]*kernel[2]+tmp[9993]*kernel[3]+tmp[9994]*kernel[4]+tmp[9995]*kernel[5];
				ans[9995]<=tmp[9894]*kernel[0]+tmp[9895]*kernel[1]+tmp[9896]*kernel[2]+tmp[9994]*kernel[3]+tmp[9995]*kernel[4]+tmp[9996]*kernel[5];
				ans[9996]<=tmp[9895]*kernel[0]+tmp[9896]*kernel[1]+tmp[9897]*kernel[2]+tmp[9995]*kernel[3]+tmp[9996]*kernel[4]+tmp[9997]*kernel[5];
				ans[9997]<=tmp[9896]*kernel[0]+tmp[9897]*kernel[1]+tmp[9898]*kernel[2]+tmp[9996]*kernel[3]+tmp[9997]*kernel[4]+tmp[9998]*kernel[5];
				ans[9998]<=tmp[9897]*kernel[0]+tmp[9898]*kernel[1]+tmp[9899]*kernel[2]+tmp[9997]*kernel[3]+tmp[9998]*kernel[4]+tmp[9999]*kernel[5];
				ans[9999]<=tmp[9898]*kernel[0]+tmp[9899]*kernel[1]+tmp[9998]*kernel[3]+tmp[9999]*kernel[4];
                state<=READY_WRITE;
            end
            else if (state == READY_WRITE)
            begin
                r_write_addr<=write_base;
                r_write_size<=read_size_input;
                r_write_data <= ans[write_cnt[15:0]];
                r_write_enable<=1;
                state<=WAIT_WRITE;
            end
            else if (state == WAIT_WRITE)
            begin
                r_finish_write<=0;
                if (write_ready == 1)
                begin
                    state<=DEAL_WRITE;
                end
            end
            else if (state == DEAL_WRITE)
            begin
                if (write_cnt + 1 < num_read)
                begin
                    r_finish_write<=1;
                    write_cnt<=write_cnt+1;
                    r_write_data<=ans[write_cnt[15:0]];
                    r_write_addr<=r_write_addr+write_size;
                    state<=WAIT_WRITE;
                end
                else
                begin
                    r_finish_write<=0;
                    r_write_enable<=0;
                    state<=SUSPEND;
                    r_done<=1;
                end
            end
			
        end
    end
endmodule